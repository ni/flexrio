`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1744 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
4PLO5jSby01Gvgd+5+tHBJCxSo22hlqaoaMkv0dklj7lMgCo6/lRhp+tw6IgOrrE
rq9AtCneWESel0+AutQVL2LtdpJ7x65bss8Qd89/9sd0E9ERwwxYyxk/vXIS9jXJ
khEvfCqzqAJxasWrwbsadk9BIB2GXbB+JyVw31OKKHrYItlJg6BK9S+/Km+aiN/J
V9EB4Md4+qHCHLBL6kgT5Qz+HBQPnuLjzdeXj7ZXkZjMwy7kg6IRc6BrfKkzP69U
jQ7rvTze5eGDLDVm7bVJDbx56+pz8dY9qaPQRbnR5im9mk4W+BLedBhffbYn9XRn
vupwhcjWI1RjpJJuKiAj89BEfTbbqObYvFg/zeoiUaiydI0CevDvENeuYIpyM8zC
zYlSDyLWKD8KYglABRpquWt/Oy2G3UzwBYTJSk1dSf4KHPQvulxzPmZIKR0oxkCu
OWc/jeDRSAM3u8HkR8IAWjTr7wRXR+9nMRIdZnE8nKwfrAQJW3AI+Y9cKCDogGG4
IGtU65F2ZyVBlWMD9U+Peo8fMk/qelq8OHtjQx0BB98bHbbr7qnK58tvunVivid1
j0NqQ+AfH8vmuFxSVXbiYUoe1qmmqm+vdjvSutLIpPtkwhlePC4hdn3HIzYoTrcW
43OPGhA2Sh9zvooI3DsEewXrSasb5RUQuTpQ3aQ8iJ7gxnDsBtDsEj5qG6AcDWQP
j7AnLUZkvA0Yi46nlCPPA5cMlVe/xkScl9XN2i9VfNH6lYTUBRl7nilEl4zsODiG
OvmjKQBRfn+axUn70q/5eVgTW5e4nHcfafUi9B3H3MY2mGnChs4Bvwu3tYMRP3DQ
gInBbvshawkvfu6z+EsPr1S2zyv2HKmmUGVtmnJ+qqc0+lxJJYoqHnuuCY76KYas
Vyam4PwCkOzG0qEHLepi6WYXBrp/K5s61eRDOeXX7KOtI9CGQuR7GCi67vSMz6Rt
shVEXTlTLfI4+wfUgMRFKjGvsngeCrAYdmKFly2Hkav1fy7Q4ez8TZ/eDfS1k5eQ
frRzroN6IUQl+/LA5pbY7Q5OiH6yZXn0B98GaSVR9dQ1C43sRPU2E+Iw/OZdCksn
QsVO892lPjI0DRLMMupvo4icleHB9QTJIQRGCiyjwXr8ESTRx3yywpksxINlqcXX
eA8aYXD2sqqThWYTO6oJ4/baSSQbd++p1UwF/+esqa8QN/m3fmpbG2gueDi/yuBC
RduqkrqUtE8N6mhInJeblj6RP2C01fe3FRfUumpQAJbAnbIqz5zg+r8Jgmz4SZ9t
QXFmmjYoptd/xELK9+9z7n18tNiewCDfOVRAiJxXhmQms6c+z+aivfLZY+yjZTQO
yv5XuMQVnmogGOBDsr9TqCgUDF98DxwDg0/2Jc23u7gG/bLA3ciHoqyas8e3i8tl
zKTxDvDPfN/HQjEbmVV8+W12lcAriXGDlFK7o0OeQoL4WwKvb3O2fht3W3IrwL1q
16zK4BuVhl3BP9RH1L0zz3e/EzEgnkzMHcZrqTkwA/DBtYfiWsUim5IpnpjyNfdl
34NlicHBqAbtBNkY0Pt5qsYyzs9ponlDQAboQJN+fFiF+xbH/JzGIlI/RhsQ4+ln
Qjkt94oBckn22KtET+YXzgxPjKN79QbZ4KH+WUaDEl+jN3sfiaw7PDZWA+Aux/CP
a3FnLcyJdCJHPIuW8wGRvQ4/PeiKeN3kngkxdblWGhLuheAjyCmjBoiNmzyCXEIw
1cH1qDsAXDXArPbOeP6tO0p3F7AAue3akA3AWQGK2B7CXaRIbkT0ZYfT38VJOz7U
uHfsuOL+5OKfVwUeE828ilprVdP21vNdS00nUgEHr1bjMm+BPsEBEoCrjU7Q7yaU
x1R9xU0+cjNCYKeCpGg38cnR1LQ9Dx4RW8w1Gkf56Kkp/Ke9+xHILiaD53VlfSyi
uvu0VqwjBDUYzJEKAyyazOO/6yj4e1/qYX2y3zqN3yIGesZVFacCsCurfqsWTqS7
qqDyJQQ7yVbixyE+vctvaRKGQ5Ko0AlbmOpmpnOdvG1EE0dFkbFaUL2jEZniFhAc
FsKMj5Q1qki7LfzS8si/hEKLHmRPzW0Ieq/UkPqjFUcG0+EDLJn74/3IGU2wBxBX
O8jqHTDcZwWLZYRLUNG3xyaJpS/wdu+30RcfCbZtliVgy/pkJJzij2NA/quJ/nJq
954zRAv43/Xf+osolwxj/Q==
`protect end_protected