`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2096 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
vdIjwSj3pLGjU3abkvXt9sn34Fp450xjyj/OGS3hfAGuYDIZ8R5aL4iueWWxImrx
xiItd7jBMinJaTYltTRWQDCCZkbZFhunHiWfFPiDGkgJqJsUQ6DJw4mHlkiPnUKt
xkGZyzE1TC0sG2eZfal88/i2qM7YEPw6gCtTBr4JoOolP2HuuJLed71q9NX0DGqp
v6JnBazBAAFbyyfxqxxfRy5T7vdySBRMsTuR4Hr99b4a7ab3pSFzLNmnEupbM+jg
Va5r+DygHsU2xvchwOPfgFq5zap2xgQVr5rznMCo1K23syJbFi/uzsAn3iUk6qYd
DTzPATTg0JWTcV04709nP5Y+xfamYuIOJ7jaSFvLreYktXTqrbQYcqQb8sVyfatU
IgsAGabJqKlKsoR6Z4YnSLlq33mRYnrD9gOsOQ04N04tYYS11Nb/wKq4QdEtlE89
3Evfe0mQ6CVAKEKBgtXT3b1ktsvgU8DDNd2ndXiAx0XzZlP+TqSslZ5e6n5PP1nW
Y6f9bq4hrVwZ+N0BwPNSBUkAV7YpBkBSEYuHNHy5cxLyzjls5HjOSFcmJVeFy/Qx
ibBV2lLvYFQd8zp63PQgf1JEx/eT6e8cBxMu22lmKVMm09Saj8Z04C3KjRJUgfHF
5fzTH2c/w9pM8jYGPk68dvvTPiDnwUfkV2tOH5D5UFLRXzpj/vk5Ahgyl0gjMgLI
6lH+OZSFsK2eiEReHhk6iD6h4GXrupsRLJooVBGv/1F2p18w3yZRvPSNfvHbJXK5
mGGAUBrnIFQYjvjJ6svurEkx/yoWrgWlS8krrDnlr8n4BewSv2t41truDV/0CmOX
TsXMeK1uNfPenQ8D8b9FCwmtGnaXNnWf/6mN91Py/ofc2bSfkOxjRMn0tXnc1p1m
AuUP4NPLv+IXecmS0tb+SVDzP4L/BH4ntUlXosK2/hrC6TQLWRs/+CfR12ft+wjX
cTaXrwBZGMK9v0Jp8RKtXOZhG5yZ3fNDh0iNr631/sAhV2Qt1BiRJ2cCnsaS14Hg
GegQwN5uz/H9yJ5SgwPFP9xFA0rrlAx03zS0C8Cs2vsyQ/ZNATOn2VdhxWn5sLhR
6LGxpZ6hKuA1LOr01HRQMqLG5/hIMM4IpTrJWpvCFCxoTqgDOYbXX5rvvh/yqAOU
NYUdQBL7ATHXgXoyDNZBnFpix6ifG+yMdgBXuuptMSNjQl6PzW78sVwkzh6fzCMh
Q6Mmc4CscsWOv2U0q02Y4UbXlbji6DnlERELfEs2maIRwKtbPoTVxnYmK6pP77lF
y+yMd4m+ObSrC+bn9RRCo1+l/a23CXRrovxSqh54M5N83adp+boB2t4rVkM3RTnQ
DlfH9Tam6Dqj/N9Ri6x5zJp9a1tp3Nqg5O4MuxZG5fKVu2r6Qp2RudmX9MO3dToj
AE+bEatLaT7JmWSSK/5jIiFX39mcrLM0LAtygAy7QiMLxSZgpMZyoCRe7W/r49so
ACTtcc5ADBcnHaK19ZNF6q8pTOI9nn/YpfTecOUVr18KGwmrArQjFIPAgj8lKGI6
FBEBW1Cdr9xDeJogFXmoBMcvdlttB7MoweM2o/VOJflfxFOT8D138/QCpz8VniZ+
6keTx4k/lAWVX0cqq4lhyC9YS97rnYwttGeQ2JGWT4SMsVu16lv82tHhcG8qs3Iy
Qqc+fdTia4oTGYRNhFHxKJUQx8HUkNOk54Kl1gX/xSMJxIQghcBZ9ZPmAzhE1Uta
kE/yIjioTR37qK5ZjPZUunwlNLRSVdb4vS0BvjKZ3uXYwu6J1T189G933fkt9iXJ
ES10LBjeTGxZ27WFHgDGdDm7kBi/GrKlgvrPmoU3v2yxCHuNkygMvb/fjPeTRe4Q
DN0YIcKZPrJX19W6zShbDi+cCMx9xyq4GFTo0iXN04s03E/3PeX3Ap6FqW0zcLXq
xKDWxk2fNVo+g/bSdWMrDegWbEBEMIpe31kX0Yc06ZxB10NCfra4tt7IXpQTzUsG
NEbaOmoI0faNWpZPL1Ym4veC1dN7nzpwNngaC81wIbMuIkFBpSZfwlCsl9n2bU11
myIl78rpVCXSgbBi4DPaJNfqFRXZFvoXKZAVV//5/43BV1Bg6HZQugcpBjLnfhU3
MPwsw0+3oHXta/CAWymCNJOL0hiDFLgCCCYAwIiffvximfb9Y+FXHMuAo8UMC6Xf
OLZ2l2l2pHw0to0UmYRPVBmXcJIhueb6JAvVgNZUdIN/HtyvAFdnqa012WAzVB7R
AsssEEMpi8lgWSstdbkYkby+MG5Wq+TPSo+ZecGA+GH8PgjO3UtYZIyHlM8YMjsK
WsFehLLZ8YlD6At5lb9JSfJQAifKE9ZEXyBgtmi2tjo/HsODo10MObVuWM5uwXvE
2xFgyNAhZxO7FyyvtLhXME1ggm33eO0VwuRNm6iAfNzRnK8sQLBtPj5Inu/Youol
XyqG5spbDvxk3Ex9AekfjxzHcQHPaydIZ0cK2gk9Xhk9GG4jdHI0FBYp7mgZO0Tg
JXeztaj/g3C2fGx1ClhTtBcWwTMDlyrbMIGwKALABButX3kYkDN/fYiBp78nZ22y
rj5Gpv94GZlKq/m+myNILjFBaHU0m+317oVLmCgKGC2kmx9ogA2lpkgveJTosy3l
E4/nKSajTg0fb0bdO6dRidnZEcu2YTu5M+inOx+hEbs=
`protect end_protected