`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1952 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
vdIjwSj3pLGjU3abkvXt9iX8JGZDwcUjli6TFJM9goUXkEE9NERFMQdVZCjtRC4W
ChYmluGzAMx6xi5uT/nqd1vtj+5x0z+lG8mIyguFTN67T/L3V7Aw7g/obau6lrKo
hLLdQw5BJtUVYgtU2W6kMUZBWlvBLdP1Yvd95am6F4FbNZgWzK90k+JvAZn7eXVr
cwcmM0EKD6Tc9hxIuHc1/SI+bF2EeOoHoHuI8dGez2gIdjjmXKwmO/5m7ksXsVBL
Cm/pvrX6pLG+DqxDdy0cFpSFufHC0+AHszCOCIq5+o3Td7+KUleWhRX5DwwUdkZc
fipVIw8ut5PayAI79jNDuLrw0Tk/tRJKACWnflaXfWCY9cSdovwFnCtqTMtqxwMz
3WsZpd8fQtZ0vYZoHoSbrtacUMMAgKgK03Ll2SHfnVxCH/ILnFW4lpTUSKllzpKH
yf8sX6wD/rVjv/diJcrKvyHmmlqeqhY5N2pF64cRQZpixPytn1CrsebjG8IqtUKe
lmQC05xH2hSbSen9S8Euc3WJWRRWpzqMPlw/ca+JzxIUg2pAh+2grHSU6OVVG2HH
sjdQj3ZHvxZiqAWgJajqkGz2n9SW3rxRCJQVZG8capPkLxugm1EIAfQFnJohI/aR
FwVU5sE2aH/r9lJ490T6/dGpLprR+KsUczBKIpljw809Ly2YpZMOv/xOQ88++khs
81cPkyPRHQVb03bhZiPIJ1Pb88WvIrF8kV3/VRSvEwy92U0aGUf0QLGqZYCizoXX
9FB2pv3kQ6Z08FrsOEcKwkP4WwSdYcSROKUu+LiT4hnGsSkLnLE/OimlARMp0TNB
DIIj9TUT3O8T/r5CwW7Ng3UiEqlauJosgTMUQ2zS6ZnkVUC7PzxkcY7wlljUYSX4
EvpqQVIOsE2DwH5fHN1EXZLyYG62GGVbV5PKqLDL/wx97Jg8uk1aQ77LMMMsfkvT
9QQTpDC/CXzYFI5kfPjwCEEOGJEuMFsOE9HNjHeykYivmAQ6PZmVirxB+dNXg90a
CQb6w8GNvu/yiP7O/iNo3nW7vd4FcrpCeELAjeyjiXolZJgFQTfjqBv1SCvNSY/X
aaNNUh8+LbY6MGnI1yOZCPPlgj9fSK4Eyp3h3WqNfYWgSu7UECrnUtscVdyxXPyi
hZgvLx9qXfHkNdJRBxwvDl5jDflEfia7rG29t7Yyg0Sx7DtIi2K2hAlJW8K9prFw
21eu1yg/NL76qBAHGAFNO2CE4LU2NRYHLNkVc7nScYEjGGehCH2L4sjFZyc4aisY
BsK2rTWO4LoyYPcM6sS9PY+rN8EDbImDDnDqDABOWy2AwQ8Zwpd4f5u8hI/5Cf6K
ce6+84XTtHxqcG8KyhgieaSxNlHfu1rXzShpRfXVAVAND67Y+7nawkWvqT+gt3/e
/rymL62mXC0DFcXVopBiEv3UmLMM2lz1eKV/+thauS4/yI9N41A4y6Wzhs4J9CgQ
/yUnKf6VGthosuJC1oARXMkQPm6SdeffdlNGHoNqngwqoGn3We3q09FiOSYgFK1X
y00HpeST9cYtFg9gnylB5Df7jwcUulzlyV7U8ErhpvsMIEVYedug7HFKyCDrecz6
GEjHu8sn80jfu7Mc8p1vfT6Zm/ytPXxoKSZz8xJKSC3ylyXHbr/Mchd1Eu/dv5XX
PaJ50SuhFJoHovAI9/WJQURWX+0zY19wBdCRBEZjzcVIFa6/D9x88uNdDFOW4lQZ
W1sWWiX3+7wuqDqqk6xDApqQQ6TpBvyzaQ+nVY8IKA1afO1CMHbXwrFLj+0JDy7K
fP9ODS8MtT59FzrH8nUuE5ibv2S0QlhJATUGQk9KMw7SOReon/jKiWTJ0LZX/l2P
+x+gQIsd9vmGBB4pI0awujbA+Umr5lQzbG1Np2q7cVu67hQbSq1mxDkhT4EbUqeQ
TyCzG1JvGVVFM+W1Cj9wIa9qNN2Tm2cBtpRvwlde46xuoLdl/tV48J+yRBEriNFg
21FJH1IBYVADX2pcnIBuKdnbPNvUHQRYFX7mQsztBBoV10SWZpY1QcAOj/aIGqDo
mgNRXRAxgd91BNwFcF8bFdTDJgUUci42g+dFG34XfyCEsXP2Bx7rksHV/br899Xr
rJiTpZEo9aepMLPKNQ81ZJA5cnYvsKSeqfcUeAu9Y+c7pCZQ/ZwH3nBcmP15peaU
hymNnJgLT7te2M2kYX3sSD3juN5oEK9YmNQEnE/EXEdb81lXNWcs8W5e8b5b6/GM
nlmDRhYt7Mfslwrx3zTtKcZ51OuhQbnNFxhFvtRwvWERwJMLpF03Lu/vuRUM6TIg
TrS7TdP8ag+NDGKOTLYn43kg6prKdbQXrWbgiyUFCveikRM53dq8Xa3dbTI9sP1T
4sEdtjbJG03xWp3aqxGZ70wA6h4unfs4rvLx8vHOSSSNFuvn90xuiP3lA2FrLF8z
noVnJn+1aQDsWWZ03qKVcO0xbnpFUnxlxFnB2HItGnQ=
`protect end_protected