`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 55056 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
S993bpJjwxtMDn0RNN54Xwzw1ki49eClITHpeOWi38ZWAhOzaZqEkODc/5/5S9oR
kXKqyf6Ck/8LXQFdMIRrF3XqyBM/xf6tn5WzjoSw9WMyY+Igi7MvKgTUiLejW5Ko
TRp3taIjsUIX4ihUOedY+Y/LQ/3IpqUi6zsGlZF5r2txp1GdnxZX1aILJRr3tBQu
jsOT/S8RwSCOx68W6p1fed6Cn/y77npzskY9kf/EGpkoq4Dnc525A2d/NS+IgQou
fzDAoXPyvJfRCFekARQB33W/uuxOEXKm79lcvlYqkYsJABVNtSgLgs5XEbB1BoSu
YCv5LFRw8t04DZnjYBZkZSlQx2dBrd/sl0wOC7lTQpjsSs4T2CE2N6UWqbvjnlZD
n40f7W58DeQ3jy2i+o2xHpKdaOHeinTXP99NCTB2cvsXs7nIs/lzbyRvretjRAYW
9d6jTVqDCO0lMoMLKfGfM9YAwrDh4BxLAUtcSSmCsj0a0j5j+76BRCaUzSU+Blhc
UqUHVtSlEwzIVOFOzMhxdkE9nHiQSJRfCdmOAV1RoiFJSQx8dhWm3Cf96KBk4sn2
2QP7LRwHfSJSDdijLBZcRI+qml4RxXh7GfBVqno0bSTJmJ84Aek4zp8NIQSgeyKv
WAD5OjhVsz2f5OJ6TWoO+FxVzq2LaZ2jxq5IpIe5fhF8mg+RGkjpW21mGikiMVyc
l2jZZ7dEEttRsKTaDCV/cGEmjbNB9az9qx1ajggQCaCggRUW/WPWJR6VR00a7Vpe
hniYmV4JJde/P4MVB2WITHJ5x5+5SelA5BCJ+42RX/nwqPgT4x68jqdMee91c7k7
rsrO89tF8KgB6ldgXCSEZXvvazBmcMAabNE101y9eXgP2OZY2dTcWTOybaAADEBJ
EXxQK7HjYOHMCBFHol5uj+nmOIK0NCFlw1VGFokyyKkyfxt/CsWaL6Hyh18amy28
CCl41xWjIy16PwyFxbsJPmRocYVJQ8McmwZO6gwrT54nS0aNSexYH4JmjVpKj5gB
xIpLnSLSbMawsRvh4Bf4CyWov4c6/p73k3NhSIv06N+Ui9XBd3vrTFsC5Z+HJemE
U4DgBtl0kfkx9dNNWJqgzg1Rpsfylncm8/1l9ASmJrlvYF01cLdOtQkYsmzPJed+
3OuqhQVVladshVNGsHDrmnrBaSdZTP4BRuqMu2e9HUXYb/Es8YkJgV3zwHnnRr9b
EkPSM441ZSjFPnHoRaVTy2YLfByDBDmfVYHLrgBTMV8x+ydLXmqZleMlpPYR1l/j
kDi5TjX5VZGTszwwiAPuoOpTKGK4pmlw1b0nUd2blCgj2AwJYX2jWvbml+Xp1JBQ
a5weqK4fl+Fw+c4oakHWpzyWkLvSPLy0Ase8XlJJsRzTE3irYr82vneo/u9evUvw
Ec6rmN1sGPGLXPvyZZgehn1KXqjj3fwTKU7JCRnFregsp4LAkLtx4+PwVybsppUW
ldDM5O3QeKJ4OIqF1jtwhAtYis6Y8ioDZf2QdSRtXmV/sf1eEqRKDWZVosOb0P3G
mwsBpa+upCl1VsiIXQP+Y72kexDWtgsEOWHjVDW363y4IJy5QjCaP/ryHUQsFV7f
9pf+XsYuXOm+8I6pKlcViSXUgBhwOkCiPWfiwwIEp1/ATSAWjmvbhRN9ZqR/FfoK
ysAKX+avbnCaXj79y9B8L5CHRvx0W+BUem5He8myiGRcumpueVONdaxYir2Sn81j
KyKFNfqCd6ztks3ldcvmsR5nBT7Prb4V96+vLX8OSfVWGPe/2VIgnl477jYloNNH
pac/o56chFX9BXSVIbSnvSOPr0mR29mbUk7Oo93+9PdELsGACrtAwoWF0CUTkOX1
oH5SrxuDy4HsdYI/f4DBfPI/BFO4lAZJFwt/kg4Sq7ysxHoEHd9lFfXQxRZp63FU
riEtBLqOBwWwhcpCNbBzrco8ReqQM4dcuBqC3fALyckIDysG2EBr8TJ3emhx06zm
VVwxHb438wzwj3pFGi/gEXt2zHpstziacRMnuC52+RgZO3ods2rYTL8PUXTZWb5/
qzgCvRdFIpX9RtrkN5cU1+70mEwXmhnjWn2yowMexZQSoehjpWi4WGa4a5DXFjAJ
CmCn/8XgnZdhxfMVofCMwLK85xM/ur91b5AtxtBhBEO3S5o9iMFBWkY5kqA62aQa
rXgb34HMOD/6/oVNE3YmoPYoPaLOnQ5NbJw9cOcNJajLIpkBI6aH2PXh0uxdyxTO
HxC0k1v2oUduM6SOdvI91anOaGKvAMwOAt4kYVsE4pASRPg+82BTDOwoFkVzgmEJ
v4R+/kugBAEfxn+/kQobChKo8g5ns52soh/pMh5BFt516LU2m4ssoqHafvYosaOv
PrOzzsWgo3CPj5H4kcZ/bkkDe3ERW8V4rUrhHK80zWWNW1SV52ot3jNv+w3niqC9
JWHp8RTdQg144MqQRgrGbp4n7sfF//QxUnt/NcjTKcspLzShb2EQ5pKtvqEek0OW
4B9EGmQKRLLJ8Jd4DsnpY3XJcQdNJsWFZS5vn/0+T0+dIEetzVSUMd1/pOq9K0Q6
FTexBxgEueGFxmSG3Cj8OSY/IMUj0s/fOUGqWrrePDnV7cuAGcBBJmWh9YUPfDZP
Yv4cFQsUu/wj83Dl/fYTIqOuIwwhhMPfpfHLtbPv6Zy/JDa17ZM5YtfL1GNDOw0G
aHvDHMACdplF/1uS21fcIqsbEc5AUCvpKRQiawA1JkM/DG1sc8PkxhbEtyln73uX
hXs15HuPrasP6BsisRxy7Dc2lLLcf6wfdPCWOp3sbSeRanJyIuVpZZC8YCE+TDPE
8KPcVpFy0a0UnIoRv7K1ErQlXN7JGjA2DFoot9keB5jtws3QqlZ/NysbOSM1REcw
qL+2vwo+O+F1/+zkB2+qTokpwmvGmP0788+ZbE3trWEw6IoWo5njlGmnu4F94i39
OXLTXULpmDsnfU82VpqvR/7Jr7F5XuXndCx47W7Hc+26Sco/tLUIQFCiF14w51bE
brp7LpryIxvgepqoV0TvdhTjgltaJWWaGmRdGUYusOF93QwZhh0oEP7SUmqDs4ax
Q5S8dpriTKOfP+EkH2qNlpWk9v7fQX88xF7+gmzjqT/zPuRA3YcR61KDmnCkpEFO
9oXZJ/v4/XHjvwPTWPKkQyHQezTWQOBqJu5HXne3DA2CcTsMFjM1/bwntzo3VOr2
MFaAd7wKo9mNfXImcdo7gH4IT5C+zETnFYygRS5pl4Gm8jZLeK0zrd1jhIDEieCd
Z/S5ZJ1uzBpwsjGC6LIZDaOb3fak6RM/r7dD6ypouLh4iGLGYnHjV+P8mt3jjwCs
mKZk3ACNNuSosoisLxCuS6cKefGNfttusOKNhM3eclw+xUDtGvKwKILaItwvNGnc
Evhcq1o/KAu/2wbLTT3aYv5yxtARyRuaoQWaT7kaTpCDBXZvxDNfu2FjOYu56bQX
6/XImKpVIJM497SYKI7PTJ9ge6SX9/z6aK/6Wg2fNM8ogISKfsusoWUeceo+6shy
NMSiveWWShcqZfsrGXGwAFvMK31LEOtyFce8zMi+9UKZYQyUQl8ibaCNkXdxUU6R
6Mw/WGZDviL/R2/ajqHhMus1r3X08Qo4DrhQcaevAg/BU1CyaG6OvUyUNvO7Xvho
YHFUj84POvA8odqflmK+mgoQA+AK6E2wBhZMT3TozCUTFM7IfKNp8KeiZi4vdkQy
ul/xt54lop+kETTiRFQ5hCFYc3evlmvDqr/pamNa7J+cwEML8UDWH7VwO3gkNItL
+8LcZy95ryWsPrPbh44w4uRt8OkHiMX5zofcLatrT+ukA9XCYZAthuEEi6CutMjQ
SGKzoST+ejKzPmFvjzbc8JybFy0cE5d0wWm5xrFxCcNgnPFgG8gl7RLZAg5vw0BN
CQMFF+fYZrUhpukl3sbjxqoG70UuXvUHFeVjioHwjgBhUHko3gQCVshgTwA97Jf9
c5ehK4WyZOBfyQEoeK2bkjgZxb/0MqOHIM9f+ZPyiknBXWlXd7nmIlawIiQMAU0P
nX32Ikzm6tqTuWJxqQBekZlv4NogJKHbsdkCDel37UgoJCld+14g4vL1HjR0ZYEx
B/YBOVh+L+O0krlg0DygUXtINCsEzc2TkNT/Pu4gvNoS2Oed+J3Xgyp9kYzD6IoW
VwG6NlGkeVNCyQPsZMvyG1iFWMK3xws2XETiTHXMRzk6rC8H4dqSfuBwv+gpDQH2
FWzqVAd+t41syfzvIaFtNCPNohr5M0MtKAATpE3I17I1n9stMo29HYhDoE/EGCCa
9hCR4oA+1NDipUrTMcH8UPGnotQVJz/c7yk17GhjCSjQgO5BEiBXhUxUdSehUXDW
FfluZco2Pl2sRa6rdCcnfHtXUg1duOBKdsqFdv5gXVUZzp27/lWiNNFRpyuQNrbH
s8OUmifkcdq9Rpm3YhMhlU7mnw6vq7cVW9YFkMtaTqVcYEi4NRxjOrdvcpq4soyp
8ClSkbn3ZommnmcDWJ8fpACVp9VhiO3Ksix+Zb1HK3hIZUGTRjG3tRNywi2yXd/K
7Nc2genNaaDH7HC93USK0d09jAK/ig6d0lzfDeIYMFMD5cZt/FFyPbN+sfs27Bnx
WX6PaQm3J2nDEmkPPtj4hxZV1OWNgrX554MLAnYapWyPRZwsksgeKBxjwzVJfEUH
FrvMJkufGA7AjHGKCh2UZ+rp8QMnQGw+qtVb5RrTBq7ISA5XI9hvly9SEcexTLau
cwT5VZpplXniDKHY0PlNRGt9YKry8oir4JVFsGv5a1xkrvCfItnNSO5wn4kEu7ku
xmvLitrzzw5IC1ZZUCyBGEjczCsLS56WPx8gPKPAl1Q1wD+Nnqd6mg2j5O0+HBov
2nJRegKEpjMDTqwOWS9/Bj0zi3xpZMlgDrMeDG3sQMHtJnBNYKOTMwOgQlj+IxkB
Jc8gc1Q+anZVhere1xpz1TC/39U2Lu6gBWWQWlHH0lWIkE0k7i0B/9Cy7dQSD5IA
x8YTUN0ev5olX3vsrSX5ilkwWwg3iuV38Co67EKlCT2Zt6myo2WjfcSAJchQ9MeJ
dTuyrzfQcpC4vnQWDO6bFfHApJdOJ3ZdHvqDAxB/H2B9qPVz83BJkX4Ez9r0CTwT
WFKCNBamqvBfTFnO+PAjBzE2GqO8G6sK4Vbble7CLrs2JXdgJFCy+hB++pSMwGxu
ifWS6HkxJkN5140DjDTFvtdM8S5ICZ1ogOH/L5uWdvXDQZD0WsIdFm0MzaTWzTkW
E1GRkC3z+ZITvZYMGvSci5O76NVIckC9R8ivT6Osbfsp1JmXJZmVE3UOMCeZqR1n
EEKoglYlJe9+EE+QZoHREGFMxqr7CDDQNhjDBUuA0Ti+/XOF4h5no6PwfixqmrA/
lNBxOF7XonXc2FltxcgLLRQmb7EVXJd2r7KdKzfB4v+G+wOu14bbyEkffITEEn92
bXX4s3QWEDuZeOaeG9QbsMq4UPyZjqN6aQSWFmkywehqD+h8VCl9ExolProqij6V
gap7mjMpw/oBOzm3q9K8I0Uzc+mJovfBhN2Ffog4ZnDQNooYmP+YGQ43GRhBf3x+
mP/sTXtXXf6sxy4Ba958534M5qHk8QXbie3IzIfU/no7HXzmc3BCGUUCQOozq2WW
j4jAtJsr9ziXZou8z/R8BqBhDuywhsBiQGTPuuV2xYVjNtacNwxPi1THWEGqv5vJ
gN5J5/HpIA0DXqNXffbwHg9cUtPFv/+o6bzAwfMJKcErDGgCSkXKBy7iLNW3iOr2
hSNnpQFMTFUc/84kMS3J1Z4kGkFIadzzOzxgYJIULgoK5VDKe53Hd8JO/rdrDLzk
xfCm2u97vZextvUtdYNBGqQY5pAX8kpragRSeXKfiYrwZeeipQBFGX5WwDIF4JJY
BrLrBfWlkoiq47tpqBwv1NCbYJLojyj26TzKdqE8UHjYRwYQ5y0SoZUVpf+DTVuq
CUnNFjau6R/L38hgRVoC2O9/nmUeQXyNOzcp/3r4GPNlexotZqXCfHJsw8ZWHqi3
1xraw2ujohWgbJVq8mvlG1RoDz8hxt5QFhHbBRtKAgX07J+sEEEzGm0MHG/TRy18
SVaz2q96K49Z3DHoTOfzV8aEhfgjY3fUUY3nohwgC1C0xinHQCI36bf0S/WjXz11
uPPZlhMPS1hPqQWAvKn3yhw2qGJjL7jmBjogb9VJVU9T2hEXUMvnmmcQMOaPgYZs
D26mC+Z6qnd47HRVMw4GjjVmnAvArixdSQdnAnRyx3TzlqgAfXVGUYcdKHvqOthz
SLbZ4UrkDFsnRhxY8QYH7mJcuT0NgPiikrn0+ckBqxeEWSbE9YFlgPoGnDySMD0P
w2t2VK487ibDDpxKeYwouWc9IBI3x2mthQFGPE6tOk+D6f/p3zYoP1gZ088vGuSD
OsHEWyamIk64fY/3FjZfigz9vnDIt7kWMIpo1kgHDwnn7HT4AZv1cn9/3rH4D54q
nZmnMe9t6dP0UXkTJBUPHFs5ajPzFI+Z1sek7g06aIrY6uykpiVoQ9XI4KtuW150
DmdsKDe7Dkfa/dtbESvPYxdmMD6StT1NZJesZ4uMlgwOoVemZ58g2RfIkoR8Dils
Fi/1VH7Ag9qJ+ssIbjOXi+uQNPaJfAt5kemDpk+t6d8NcWV+HXja/DshHM0xSGBK
BUZB2Lx5JB2DdfCxVeuiMUEzmPMn5lxeVK4Pz9v/krEmXN4JkL2qn+9RZWxLk06y
RKgUKiD3VlSWNFaluZ3tZbLHdQb1wuzkwq+zm2OIDPlUpVVO6ZH1WUGfQ6UMMr5O
rZnkY044sYErdV0Huam2t66zHf9X25gFIwCPRVHlFzb3Gu2z1O/zqi9xB2zhGhUQ
3cyu+GgNAF9+vNRKyEgWYdz/1s1ktdWRM/Vcm99xI1EVNAL4phqoJQRmDPdLUii6
cXyd4M/DAEdgdV6RYL7iWz0bagIt63tS6WjEvYo6AT1Pbtz9kwJZUckf8lQOibIF
L/GOfIUDpm4NTqQmlDfgcqGW/vgfVMC8HZ3oBkTJT21iHXQ1dyBm2gv8gwK7op1M
5IsBOrOiPwFYS6JxziH1f5LHi6YGrYlvmTgV+rc6ZODsUHSaNtwduj5S0wHkYO32
aN5wLRlOFRgxUz4E2TEHGOUEkyH6KNwvuy4OqWLPTJSQze956kesj3aWT/mghH5G
xImk66XcFsjLhSdQDnT+Bnc+oNft3eC6JIE7BCyz5XfhWU/kT4nob3NW7naLhsSM
bknjJrlDasTg7HnvhQG6cmwNPzpNqtamtbFlxEqBVi8sA/t0zfY2WOuQGd4LAntP
sZCq8WoPpiM9TzznZ/4OqMbXhkwwvGFdoGWGi5eUeitvoNlGfz/R62KeiH2CWVH5
eC/cv12rUsWnPSJQKUhl52Lm2pBDPdxxAAriYZkANiOUqA7YQMCb0dgfKO3AMdfk
XifXcI5UOC62/0HMPjoun4GsYTJJgWP+zRaQ0aPnAPs+XMBOhJJualLhcl+ejMFC
U3o+x3s9aqsX+vZAkC7/ks+0bBV0sJLh54nojJhmB6RxF7WrDO5scuepSYGeYC0Y
PmlfCsH0H7HRXRfZh8VrIqzryCCsStHHwMfHnLOicXQGoNgFbspFQUbqExdnKDc4
BiJ5quK/S7emkneDcOR/TNFlc1e3d9QRTmwaX7531uDrxriXQ5Wx50DQ7QobaGTl
sZQrEBZBI68eMdm/IozjoLKtb5eJFiwo5Z/zwgf7dkhWb9xlwtBxsOIXTn/ONioj
/n6pQCA5II7VwgT1WEjBjkZz7odH2b3J0wfSMVbS8MNYzqFwLlrIVqHfo1ormc33
1KtbIZHP8q6sdAim77NXgE6h41PtHLxD+hg6ibE9lcxWijSODSdF1p/wEPfX+zAg
1Xe2EAlRXt0BWJirstDT57aZ1VJi45O4yEjk9Z7cri2ZVjJBbe5/eq9zL7GhDnkz
UXdeoqImVGlg0CX+jU+cL9lfMrlJpmPcpbn1wCP9G2PJVs6ovzE+2mhjqlJvD/2x
t/eUXxbEUuW913Q460J8G2mpEg8V2KtyOK9X9jP/DHsydeBtzhdsYV5ejiirpl93
u99UT7J4AL7gh7MYcP8PqXqYRtVfK9fFbutJFM3qAAya+BknSwnhpSiMrVwqaeEX
LzdAm/Lx/FnUoeJXuzEV3DkwhxQi6uQknHYXK/N++ZAY0mWDWJtrzHikAznE+m3j
/beBOpfydqQroTfaCPec+oxRtpDMGsZC2Aoo5wzB8uhU9k7cFwohH65LhRgCTK/B
TEoWFOr9eRv57m/xAx6AdLbHYgl8MjzJK3gBDyDZieJXco9wfw2lggf9J8BHLUM0
nnON5UDxcua13ZDD8tjtFHZ19XEKssJbBk2S+kjI9yWcOWipQxJTovRneH5+uLUK
h2lsAywQcpU8q5FZmu2wrYE/FZS4BkB/Yx2WqtzLfKNFI/bgkdo0Cvc9Xvbx+GbO
BWr74+E6rfueIuRaNl0EGy4ZpwDO8gp4//odi99NzFRV4rEYz/44pWrcWpcxeRr6
M17BjWDF2Lb0WzSxaC/HLYicPmqfzZw+RiNpfot0nteS1wSyNAkRr0dB7v0kwZ35
maieRuoUFArcteVXYJ9oYq818L6f8ahxXus2grU3uLdNhcHMqZMOJkYjfsspAqIO
tOeLOPeQZL+U3VGiG34SAiF81wGKFtjOm+nMsH6qhIruP5kL6g2fZEJesSXwS+Ch
JQfwAdhYOmn0hqrHHHdk3/NYlALEMx8xtEKXfwLqzLHc02Y5QpXkW1cyOP966cgT
C3i8prksdQHsgq5uDs7zfmPUyuMPAJawgfIBBBot1/uxQDlvFhq3G3n62w/LO65N
nkgLjdWVZlkEZnQ4R553WiZCP+PSroQRPGn1XxQfosAA24QIgO1UAu6S7U1mfdbg
KVFNNnbDNlKL/9RwdvIp5EjKRh3jUHHUXpJKA43q9koP3SNCR6xPPFCdbK2dBCLx
IALZ40j5MvbR7IzvnBH6I+0nbAh8wYIUo2GhCqjBpKG+2yuN++htL9DIFrTmxLsv
8JCThS6YV94mCWaMLVLFDu8LyxD5WqI7tOJHDWl//3ho+jZgTpgm+ZoCBkyJ2dUP
gnpFtx4P+T4pQj3vREZ9anIV1eMcJ0Vvk18mUSThlhoMwT22R9VoNAFrYonopU7s
MflCfJFHLU4QDUEBGlG17fQKu3+sCjhRdAx73iIdJy/qrR6AZDR6o65hMoYFeQ7r
h5B6YMLab1dmFhPtstNWAvDsfkhJpCz2bQ/+G3dGCOTq7jHsaqDex0DEqKmiyfDS
NlwYlu44CWjd8H0TqrY8YI0/pudij/5dMX9QKAf28YyeX5abVPCFrrGYkFcrI7yV
xsuQGJuWgG6D8U6wLdPqZVOaq5ZIk7AJ0dBfABlG1SfSQNLVdnpWyutdXtT0L1qi
Xw7gX/HNhXi0K5WU8Fdm7q97Q+Nz65vHcRTHgKWBkgmdT9e5LZlJyiKsO2z73q9o
UOADy6anIKOJm3IM8fy+niJ8c2FBNYLmAG5cAGFPizqbV2upbbQaj+nNOuZjUX4C
lFkXunFCEdO5tUZ2v4jdQfFXo7fCwDKmJ739WwYOaGeVn9g/YoQF+QjFcclw6ltZ
iR9ckYThn4GrVSmjCYqNTfING12o7U4I1SJMlgx1K85HYyZs59HO5d4VuyxBoLLA
qMLw5n84dsZ0pe8299CZuxKm3ECNn7phOtXyYG12g3khbGbgLivC7Jhx0Z91GizU
OSi5iErJ27ybXc1sgY7KGJ2gJd/qlagLH9VbG+Mvu0Dqd/MKy1sGIXJP5QBISERt
sTQDa2tmnq+yJ6aJB8Fz5YJ4KVKqewtAJSaikkLH6UARoenLnKY2Akx0e7Y0I7yD
4oWHsXk0VJUZmpViknwMGWtJtlRyj9QYSBewjjUe50D5w/XBWu60Jo2NB1eMpt7E
zr4FTgZoGUI9JmQ2DAIqHN+NPw4BdbAyq1wuD6YcG8mo6yVPRAuT17LDQcYlZ2LC
ukoTqt94l2GajZJoGKmwj3Z+38klMRcf3jjxu8kjlxCpCL4HonFiXvoXRbev5BtO
BcOxjDggJ6mW7yJ2Sl8SbNkCcq7yM/AYCvz+Ytfm3Rcq0Cpv+WVyGvUAT85c1+gm
3BirxwKE89dfK4fkBpvJzMCT+ILEuRGsFrudZcUfz/6pie4j2HVa0GgxYlSQom4n
20PmVR6/jH61x7By1uzWQnBNznokqLG9XhiOuQ45fT+2LHHxHbmsZqPIw8yhbONr
ElrDAPc+kMA74xdvqPQG8905t5RndtR94pqROtBJSErG00wl18d+DTqoFKpoZMZo
JoAbd40nxBFRvXJ623yq30h2lRaWxJE1dFydaT0ernlqAFe5wB6+Vb6rXdQe7f9X
sQwDigZmTLqqEiwIw9gRgMHa5t8fIyWcCxb7cyX4OSvvUSn1lPvemDMZ9bpOXZk0
9znDsg4wayBqj4ee9aFC3jWBkM5d2l1Sasdlq6GQNn/e1DW1uLzf++Wt6J9NcQLt
Aj2UcI1BNrHwtADete5Z8fg/YoMeISCWkSJk9EHYZCBhlm1XBc2YFsIYBvwwf69D
MiJvxTbWJ5ZlMs9r2ZL4Jn5n+BRlAWJoFXm+Rp0PFDvIQrKM0Gb5jbP5EnAGhqlR
ZQ0U7L+/FA/97i4WCBgarmMSZQCjUPHVCP6tOUEsPQ/GnVrsNqaKK/gkZE4GhR27
MbqQ7sqiKV2MjkTH+vrYQWSoNMEe+uPW2QxdKCzpx+Cif35WUmQG//2+3B/JY03/
B05hZdvPDP4uBuyxYOeK4PYqLSbJ9e+ZEqK6Re4ADAClWFbd6ioSpZdqxeOFFPIi
cdKNUQDx8S7txB9TVlaJxqJVkDfEk+vMg7ZDlohs1lO4/pzW9Gk9BEItdscZzJdc
KwQnVpjbONjpjn/KsPzyig9Du5X0k4YJHo9+jlYjImmyWlqLqpIEyExcEujkqPXm
g+wWhAVGHf3J9P6/PB/tNwvoxuZzFxdK5CwrfVQDLK5YxcnmaRyt5cb1IfJfygnO
F8wANK4O3SvSmuR2uVU8P9w1rxUZIq7Yxhaz/OqXB7izJEFc7M2ml1MOvk7z9AcA
Apnly5IQGReNKA3UQlMlaQWfiuGdbrw8aHXVK+eAbvHr6lrp5IgcHd5ibHxvt7So
kqoLhCcfM3jkloE76ZfBUOjzZAOqp7YmVc+H+EguPEuAy0rGQSXbx46zoompgpQB
7Ht+FSLUU89+z1BTTvKclE1Ys6lYyaPqEm5KMCEt5/djtbDHyFeGvSJc8GO1ca+2
rnI2JVNnRoRXrltGrutwz1vVsQEiVrPP1Pc+btTKbMILxYAiJd8QWzPEZJXGEH/P
CigOWeHrJ+R2h15oFEN+tN/vo1MKFHgQ/3CLSpUaSztL7S6qfTFhZovbwV3SJrcG
9qvJRENfEm1FjNnMP/vw87k6or406L0jwsCJ8FUJ9SEwRH/PgRHf2rM3gFTIgxkq
saUHXViZyJX9YfB7dgWd257+VLkV/XkLZca/qY4mDQ1cL7QRShVDxiUBRKJxqqQo
54+6V8y/g8W0DmcO49CVdiIlDKaMDbUPEJCwunLB38cVcr/VfcHxsWiMPhg7sQN4
jRx2nlzmaxB6sO5S8rvkMepEzzeU9QmO+O+h/9vfS8F4QEXcNYOj93UVpSasyu45
XU77/8vTzl6ZQmQ7wGyOI7L8/rq7yYpjgcKkkUKAusTJSOrfisXPPUDq75lhAlhb
ukeDCJR1JZvyuIM2E2vrBsoqrl4vY1qCKTCn3IQPuvOPu1bUBqBvtxv9iDbw1gV/
1IWzHsQ8Qjm+QOVr30y7L6hmVwPiA+qhKFh5Q/QcgUcK1jsfN3/mLrsqiZErTGKq
6jByViCCiaUPbFIvVY6aR6IBy+ivGvZlfo70m7fBffS6UZwvvkddxc74tfYpNP4/
+LGhKT9G8zYAsHy20vcgT7v1xDkDbNp4i5p7kkPRCMho91qitn6ACCIW7Vy+KRmI
uqiF4kgizkQhMakRVqPqPBt63KhMPzzasz0xJagZKHQZloz7fldb5sl69VTmyf+7
3VymrmI9xavgeZLv25gx1G5qygHsWWsG3Er3oQ1VfHi7qKYckDwKgIO+XNTBAKCO
/RVTg3DmFLgso2QbXzzzNJ6rkO55EPlx6+UT9QyG8dWnibjfkDehW8Vz3vTqEmMY
4Z85rkPjSDYkPXItAbzmrVDGjSnfcZDfu2qtrkwztwyIhDi+qV9IfrKIz7y7BIIB
OUUE9mAsvRooW2n9yjNNvdChii8hyNn/YKreXlRsYdrxTWauVIyJxCCpnGXJe8Kj
NQTRhuUKur5uEQxYyp9zyOn/kHoQsY4VixCDVzvDnuUWgBcHeqfKBRK5XpknjG2l
7owWF5o5oy+Qqsb8/rmsFNvRTL+XWLT5d8Xf8wOMwhbS1EaDWokZlh7G/S/0mqx5
qBgG3ajoRwWn9UASaQAbVYVI6PxMdvMk3bnR6QCQ/Od6NZr8cFG9u4suKKnyegC8
1SN/8cHUQdjQ/PNVfUNo5p1KmhySZx8iH0ooOXp1A1/Z9a/eHt3222tB1i7mNfEN
59RhOhas52CZWKBt4uFH1otaXeS3+jCmX1eLQ7U/iRF4aODeyBSiP8ySty13AlK9
FGv/RFPqoNEFE8ZOHV608iU08qAhuC+cV7dkTkworEVZQRIOTSdyl3dHMpsUqu0q
ddjac4F/pMFmRgKlL2K2g8NyoIfcBRGqTuXnZ1oxEEGVFs2C76SaOyTDZiid6DC9
wDWV2pVS68Dr7cpsMU+n2oCdud26sg3ywins66TxJKk7O1PDo10u3Id1EuuQgKmr
xAUdE2izXC85+2QC7jtcFxD/0+DzO9MrU/q6+UXlOlH8XTNghiW3IAE1v0+rLqkF
UFAvmuOF2KNggwlZ5XpMIhxpvEnCTAG3Z/CGVQOaXsKL7YnZdSC8zZlnlGjASQKP
E7Jvw5h9Y2Cq1UWHUDeAV7h+ZGvDlH8ukzhOS2n7SZ3rq+sFqMeLD9eNj4GyoUKz
PGF9cFyvRvFMIiukTrEyayOZ8O5ClwxYoHDxnceW/dXghu3zhxBOU0MzmHkJGHSp
BktjGSqBuch3ZbLRHnPHCklbohb5qYx39igO/ZoBzMoCa4xDLku+iiSRyu6ScP99
66xAHlnx99tc6phAE2+ByoLxZNF6KBB2jk8YdkQ9qn4wazzJ8qpachrkzWiM+9z1
eh3L0Ss6X8bhSHvkuCJjOmpfCp7RxgLR9OeUj40jDjK/wKmbkJ3wzuowmqtOJXzF
tv/kYicwyAb7ymYoiXJysOrwbfeXwBJXTfzyJREyl0dQng5hqMKeCUvX+FfZyu9P
+OIOej1ANVUb0kjU/LA6Ovmlo7QjbbNQ6ShH2TRlDOvjufofJ8OinPwOFLialhjv
cZ8KXpGkWxLNT9bjAWlfl5Z3ntE8OzW6VaanoMDJUzd84h1uXtiqRwpDJBrgsi9S
WDJndnqlgXMV1GBXL58Cvpt4Zmbk33mOnK2crkcNcWuiahnHgZAkRSnTNYf6zypB
pZKUzAWEhr6JYT1eYm9ZkJeZCi2AUWQtskkvo5rnKHyLBQE3Zm1MaOfEB78Az+O4
xdqknvPNvy67Y5V/isBiSyLz/xUzt8VYOipKQUCSoJebMeeHavpwOyx+fpphVaaL
yqTAAFUkC+Eznt4rQUU9guKQR2/RhJe6nZxZHDfxKpifGqBOzoh512aP6xzs1Vk+
hLqi37jH/cUwGKQUcQ147y7g9YGDyaVdbstaIkw4HlzntEZbcbmQ1IqmJAvQrLpB
zgkj/sgflpduOsWQPUiupKSdmOoKSC5h3VLmDyYTBCpm3EWpttFDo35w1gTXughD
iOznJPIADs4kbErWq0UsnLe5eavYdeq3wK6PZSByu31jAEHsPkVcXl1bUuStU0ym
5pPuqEh/eRH76R60WzvNH4xRg6yTk3vPuGYqb1mh/DDjyIzdoGEHDCRpPYk5NrqI
15C8p6sAI1yLuAmqmRUMsC4NQrRSDr2DH2E4JyrMxLit02NVDfuO8alE5DzCRprZ
Sbsw8q8QZpK1CmNOXufZh6cpL/J/0aQwd60jWxq8Jx86OyuC3UTidiPzUIZ/vDAk
Wml+LRBCy/FX6L5ANukSWIZkIidxcrw9Z0pMinI3udpWcjdsZSupDuy2r/BTDT+7
jITdlvrGnrZVsYnsMUTTstsxVCcNlQzl2kqy3emq8wSClJ28bY1c9ryPqKXRJynS
UgAIr2jxcjxGGEt4oCAXD3LJAbKuKhx+/6a1VWkYUX0zc490WRD+YpU/UPUnUXcp
KyI0u24GiSmQRwirQ9adS6rNUjsF26RQN62aUrSX2Kjo8GNvUGv4zGcrUsxhUBGL
i5jKsNQoxoPg/r7G/hgAADf67VVSpLOe6vzmLVHyJ2QL9PcngWKKSRggCdpCTkoR
PfHNhYt8LHWpy9mev/lUuEHCPG+R/VvXiGFa68/3eg8mGuaPoXT/l528QNViartq
Zh1RXl8ZZetwXRBGEPv/BVdczDHAGgT1vrbkJ6i7ilUo8UCsa0hO6DSh/QltFuGo
eEiyH9/Y15DYDITiP9l/czRrRTybSgOoFAf/im8DU2/zMryls+gSISIvZ7dVOgKn
wd2umTfs7JiJJNVSLcpfOH8h4FYQgVWnCuzkihSNZRzYFV7VWYBNsQrZiyjLigoL
+4FjY/zI52MPZNPq/2ofBMrviNDDbyhTVsJVSTei3z2aDmdjcO779Mv2+J7MAhQC
EiiOJLzHFsXBZn3wIeH6Y9LcJsMiSB35MddGciL0WQHHKM1kimcYc2Rm8N1y4liM
6c/k3Dr5iHhUUGZryB/F2yfR88A6536on0+g8ClnZa7HaCWyrZsPioptgiJkTKFd
EG9JduAH0oT0vipnnJZsrtQ5LdmE7CO5xHp8X5cpY00rCHT0rllAn5agfE6DN3V3
1x1brOvr4722E7MmZTz2uKDl2+xmPi3xYNp6nSdVJT6g9UXdbQ0tweOp/vZPyRaB
WOY5nrITq0mzEBN7r2pmXgL8nVKZxHGYFaCe6hh/99UueuVAxeAq1xIO/GSE8j9J
TKTJkXGorGaQWBE9FKs/Dx2sgA+tjEiNeVDbOdiebTHxUnaqw7noD1cfb1DCgq7g
z/nloBiaUfna4N/BjsaC++CyPlq6zE3vqguXPhKAiPVAXboBwSTbiGf73HdHdRiO
Uxx9yMLLJ0NQiO7e6H9fMfQsel0h6UBWi1trhCYAvjkU7mh4TCB2W1kscoP8fImP
zarbEgrIWQpoztZrYrPQxlKonrh9Btb8OW80za9RXC+RvkvKklyYLdoBRYa6iuqj
/tkG/hU2GByiYjjVQfZv//pnYrOo7F0ND1mZJnkXGLr3WmnbIu+kHKBXWATPk6b7
gXwYr78/62z3dEjjeNmGJ66Rr1fiyG53HFfcRakJXYfOKT/2q/JnQimYAqs3oOno
tBrw4/6y2n09ewK2wvsisp79Lo7bgHHirnb7zWUq/fsPmfPpeb2O0e7/RP0RXABi
HhN4Se0lauiA4CX8mtqsuRHZjEwKbFemfkR4V+JplEOu9O5zVQZW5kIizcike4jR
ESt+SFgCTi1uKEjxDFZsjm3U5VJHh0VEsThg7tyaMnOOQClLmd8jFuPbSjGxrtiF
rwbLpftyi1owJk4UO5LSE1RdsYiZispiMLsvaAp3N68pB8aw4kBCBuUrc7MhmqBb
WB8agMgovtIAgok5uj/Z1xB3apil6s0ljxD29XXmUfdY0Bd/AnuJpLzWhsF/mexD
tWeGS/cRptoc/vjr+2AUPk6KuIszxu7wmrPSG3XzLunxOuWYio0B49qcJ9O2s8GJ
TaL2G737ezUcRE4Ifdzrrikj8j6BXAW4jZMeX/z7gw0BiWBxlnr6DdaFaESWlwb7
tb8xdBAQ8PNsllqrwsRDOqNQC2HEJdG2Bl9CJ3d+Ns6KJlMcLF6yaQLODPfOckOv
w3qrwmopMAgXqlIbVzF+ntAX/9GdI1M//0hMVu3PhjsbP3BGp6sRYEGj4BQy5Wzd
p7dRXLyQh/qahM1KCMwWWsPfVf/Z7pUdQkAB6S89D1jh9n1prWnfQk+aVu4ZugUu
+5fhkzHO7Sc72Ng87WffVPfoMQo+RYqERdjFjAzSeUEAK6ZdNooBJTECbbka9TNV
ZPJleqjLs1B2UPqBijDNWxWSZ8Z4LtI1Yr7SOecMk6O6YxUxj2UE/HKvjA3qqZ9I
K0hgCsIKgdT5rpZYUkjqXsPVcIoxdMwbrISTt61J7hXLAuzAuTVyJ2yi4ddTFAlN
kf0x+o9EPZB2k8U7rNh7Ca1N0qyjG3aXAoFIIm6arHjFSRmkY7rEIMG0U8+BdDmA
L37s1X+n0dJbt4ZS6xCt9HHZHf/KijRm1GlejGn7Zl9HwNjZGSj7qCT8rVKvEEGd
fE4yauNGQMJ9SiulYlG/Nyio0JLLeAdoNcwHZ5cnlCnle4db7UsztQlJlUw31n1X
kDzUsge0Oph+tqNa/8eZymgsqQ/0dK8bR96cVYIqy6bcuj4bytx064KGwTUuwbYw
L79D7PYPvOdUI0rBK8Uz4Q3CPtpNZQsoICaAteOMzOsk/rHu3lm8HBUzW4f98Q3d
8TZ40xvBH5+2dWWEQFs3jzY8hs02i+v6N/Hg763BZTDqYpSzggghe5BtuLjfvnDG
KBpjWcAV1N8f3kL2ZnbH7T9tqdbtMMLrkfZBj1pjHQyLkT9I3sVF4JpExHAAkSpd
rDz/4CxPVPjdaWTRGtf/sHH+Qw1jL8VGGbO2ZzhUQtn88fihg16jLjHZR9tmSUbQ
scfsO24NJkjmvjKFmc3KJz2WLklWM0Dy0lPwxF0Idkd5OH74h4TZiNzbLN3yYcsL
AbwTlL47JCwqls0vjujV7L3YzBPt3o9N3g6vgyGwzNu1hV/gIhsJAD6NPzo+zSNC
jy4SlQ/rbC4GYmME+qgmSdjAe5i42MDB+ikoNBwW56UtGYaQgtjXmf3iFpa8JEzP
BhtcZzlS3MU/Or5bujeHGQzlQsTipFfhVa31Dw2QsUB9vRrGVDRsxp/eGVeBkFoW
AXgQPzqC96FHOg9G0fd9No2GRM5OkSWHksRWLdeMYJWIYvQtXL3pC1AtIIvJVQHh
pbt8NHoESR55HxeUFQcO3czw8Wsyn4SSw0j9COMrxHnyA4P4LIVkyFGVGvfWFLEw
yBZDd+wquJCb4xRQbd1syYEzR9KVLrsEGHr3mesL/uOM8rdLRdddMhESAHkrPgtU
p1r3sdhSMN8UcFiV9fQDSQfxdXZzKqL4xm68ck8g1QkokL8oS6r1qOrw4zzta9GC
bEX26/r7hKf/7rrW+eXEubiZoYXXFQDwE3Cw6B7leOBucMf/i3uj2BcQvg5u1eyI
Dvmtqz8+/agcjmhU7lQyoLUSnU2pNSRoOSIviFqaM5Z4Hpmi/Z5qbwAjiOyNrsbP
80oHgU64exFmZ8DSgzimBSc+ZpjB9zYKoz4cYE7eE7mepuQztsFCfzvRFalyuCAM
ftM2O9A0lgEpv4Eez3EP6e2tkImsVyx/eNT/4Z3vT5cXyXii7WCv5x4lnxqXnbQx
3cZAtNRvNrYOgeMuHJQ7i4dMDCDiPjNVcNZm1wnZ1uhEYZD/mVqPyp3X4Nls+XNc
jHoD0s1CiKzdkJDENJS0dNthk7DgroEmXIaxSyNuEMgBHOcBZmsWH2CuoqBBtnSF
TnRO+fnohjQsqR391djbgHofJV1d4ej+D9QNAfHwZwbnmUPmUHlc1Ac5jPIv7bcX
93bfnJEUYgA6TXdgmb2ZM6XoHEYwVE9oLo5kntAUUkmOWvzjR7uR7bpdAZDjmwg2
c0MY7aUztEPmRYizjhe4uDcpqp5hsLfxL5DyiECWetYjMHW60U3pRFqHyAdY6hIQ
V/FSD/jrwbiBWXX1J6UNKd+M8Qyy0rDVf49kRi1QlpZyzaycn0MIxXAMY/qFhIM0
O+zzONqNV9eOzvBAPQ/WnUOD/LNtzwrSd6BxdIUov34y2mwoc8kp40BfRwsbpbFQ
lNGNsc7SvwWQsziLOvuQHZqqj6/b8TCfoeBizJKhLEP7OOUHOw4hBdzcphXMZ3wJ
NaySv/MP9/KWhWfNqDIfK5XV2civsHlgIzI3yqkYYJHOsga8kFDAR6BGZvqvQQa+
rBJ3Ez/UsLCvEBHZXDfhhmFORirQL0S0l4Nh5qW2Ixqt7LCLouN8KU9/IlcEeCOL
2b5AVmPP+E6e/UH4uoUU3LUFlGIKR+HHskq/OnZYsyCjcV0vpK0EL8NJRP7inhPu
0euJ4C5qDEz99VPA9GKGC9d6SjuNGE1woaDpgx+PmhjXbYO6qQaL17foq55GAoiR
4FZbqe+RFJ57etKFtxZvHdHv9oV1JEO56wdWjMY0V3yG3NLfo3v1isdePRvsZnEZ
hsQiotvV7N7hyogRvnxoOKw8XMiMe4A9pYqJ4pqp3NTAWBMlhw1up5F2qVBDbsp2
hgHmWx/CZ0wPOKIU0wW4finesdj+v6XGczqMW8Cf6rQBD1HTkb+E5sJBLDwPOyHP
RdB9ECp6b4L9xypc0M/kQjIb6b6DFbP340D63aFevQ5ZIoFilWjGR3YwSENyVdCs
ba78ftnu/wMpKa+OyVKauZjnMTbdQxhxp5xn6dybvBNq0Mq76OSXYFu6YgxHyz5i
XIQHMZFouGVmyGaZ0rhfiBBaMiYBcwzoCiFDKQRxflfrRC/w4J3aYUj6ooeTtbW1
XXo9nCoKMAY7dXFnf0xaDnnZR5DwtaZywyFrwwc+G/WK6CEqpuJ0MalV0ItGkWR0
Dr6cCyaF6owbJUG84mP9KVg+Pe7oHrEDquxPBzJb9kw+egydmWxINaYvYjpYTXej
Lbd2drtRS3Pt3Hz+ZizNZKbDrHMPzLesWnJ6Mk8zUtnohh6dET1xynulFw9SKm2b
I82PR6YrLCav3HGLrAPYhXy4obP1lcMbgmq+ma7YaZ0M1p6RszeVrXt9AMW3GVm8
CLtaSxckeAvTml88nK+XXmBATLt8oUNeG9AxLhIagm+x6JZymcE7WU9rTwcDTTTp
OwhDELtxMpM7Ltf3UdmBkX3g00H1MAK7xMkwbqwiMYETOjjBTo1PMF98TWU6TTjx
kRwYmDy/vnGprNhx1oYPMK+xJ8pBkM75gm6eJfJyuNwNt8TWHJm9K802QlJ2RT+s
fp0FXCwTvsq5zPGeeZtzIo+aiu/ax1fT+Q7HgY5DeINUYn/l2ZSLgb922fkAx9+w
oee/8jVWOjvTh6EqM03cFhDodz5gi7Hf4BwaXk0JbsU4BidJ+OMwg12p2bTOMCLo
0LjHAEU0vFfeYfbE9Ce5JydKeB+lAHtvAP8/3jHMYYYnDVTQvdCUM7SDZjPg/gHr
DPfbCwKU6AXjw0WMkiW/RLxyacfkg+gSH2NhCgQ9By/bZkf14IOBoCfdFp0zKSL/
f+caWccnJ9oKhwpiBx4LMcTp+E73afRnd1zAF9A+Be2IHkCzDCjPo4PCaPGaMIol
1P1w8eHNrmT9bJDLWfLI6K4/aMvcuXkfVoxiKwS3Z1I5I+8LQIZESd+iRPwaMqIK
nBnPAnw4NYTc1OFqcUu/pC4EZk+JTkRHQ12uvRfIuY5WJYJebJu9O8DKsJMEhNua
CD/MdH0TSejSHqMkVIhm5KMfQZ7JYcPVMCsbZgv7NRWZIwdkzzPFPak0zJT4mvGs
iWHGYR00fYPUdXAGP0mJ5YCutN7IIL+MXCbNsWCgzmDiHaZUSVbwneG+PX8BWibW
89DklUDOpmpMWr/oHwtR6jITCLhjfDxYyByhhc++69mNUFxSgLMxAfZkwalmOC/U
yYHEJFiXyTfV4D6Wli2SiUos90ZaWRKpBnhlFloOvMpR2OIuXfOvYiV6JElg9Oic
T5iqHvrno1252XlOK9cp1hwRbxO1gjoOjFhQs4WWi2sCpfBCLpiWEalhuOirK538
w77kSKvxJBZE5g3QRSrQXavl3n+1mjRUSdYRMIlMhs1+7o2ntY7iiU+81MkcvnTa
7UXxRFJKXF5wbjgzuA3a7jyf4rvl21/A2KMoieagg/biHvoYqbKXOStxgDOCtHgB
pLVzLU+FEknpFUn6M2nAXjFlJEFwh1jP4UvPViCHLtzK6UcxGAU4/KSI/jIYsjk0
mg4DCfDG/cjCrWyChYWlHlVhnrQIPl45N6mTc21OaAOBldyy21vapEaADeP1Y69q
M7PSW4bxUt0+LQz4OYnT5b9bbAm1eXXgeN3CEN/VkLSLR+R1HRKrdI1+4Kpuj+zt
PlEG9deICnCe+o/yT4J4ld1XWSv7gzv4z4IX5FvQuV0peoANzrmUJOl1uvinFq98
sPrzeKUuA88tZXZCcRL9d6dtEsbjRiainwLFyGHJXW4LFD8IoPGzRDWIG70MoAsU
r+XU4Q4lrQZqMcL1LYJeIz1E2ejnlCZ2lW8ZTr1CoTaePDxeZzAgOWC+M63ybuvj
ynaNmrDo4aA1QbZO8i2jDH3V7A3WEd0EXYymZ612ImxX8zmmgH5ABOLv+eaylsBs
66T4BOSO5LxF/jcRRWMrMhxYNVbIqli1W8p3TpO+CHV5oRYFbAzetOSYC3xz6g9D
lNCBA7mLl+BRaLgiDDYMbCRDnks7DXj+dQ6l3gKEdUK2gtA+sMPqdGFxdW/6Oebb
UfeMPVzxYjcBXvrY6ar/O6jmhCfnuOM1e/FoP0+SIUi48BDBnGT1Qb6KdCVUx1ck
VMA9R+boPZYijG4n2MbQYtJ9zsVFX7bWXxv1ZpyRB3NmFqPY0E6M+vpSz/DdO0v7
/TyHmMh3K8av7WVBDy1F5iuprRaL5MbUJF4upr9SPZIvuN9eFwsAXrh65RhVF8yF
T+/beeL0a9y2Og2UKrWsrFhUmH+9Iowq+MvXvNOa9kluzUjvyZrAcDeAHEuM+5II
a9VvaiJdDht32mWtDCwVgknzG9+TB61XQGRUMpxdC73AbGHVVFZ+R+dSH/WGd32+
fBtBhHgDWeeT/maLKonm+f452dtEP/PVU115qmerdpcaXlYoWm3GiI1Ks/kZPETC
m1l7D5Pg45spCs8RYxKAtkPhKKzUIqzS2C9hb1IJ1t+NfFQgC2hQG6I8hXHJ+KsB
tSIeIgohFnQP7tZ4qSEtQ1SaLm0H73yYPTi2UA2QdUPevs3Jeu8oyogW/4N2uVzj
SA+6sLt9TZic9QG7d4kJ++Qsav+u0UCdoAtX+IvB78Z+8MovrxU6wsgcWwIFYlfl
MGSzlVUkXCw3PrCWAGhn7dHD/b9Wg6L+CU4ShI9KfcaMIrQH8Lqp3GiiYL6RHn8q
7AQla0t4lMB9SCC/khY1fhl20vnwcYJ4f9FuPbIKCzuPierfkEUvWrZw1XPWhQll
f2Tq/H8o7e/8QcUy5XdN57RGSPR9vx+6Z+W5JaVuFBUEx6A/co1OfS/tGwm8YbgL
aFme7fvsAhAJHn+sCs8C+Ns+I/pSD3ej8drKbv2iyuavjxPc4P0RXX5vjfKwkWWu
jPKk+j46/WbsFNSnHc5udA2dFp406cQgArqTdS4/QktFgwX1fDUtBS5k1IUIXT27
HcxNjc99AiT0JlIwF5B5bdv7YTBBlsB8Yd/c5CXxPM084DGhGuNHNijG64qBYCwH
bfO3PZN/Lgv/2ICuXXdw/r4LEld898m2KeP0TjYcRJ8uBMVp648Hb3KmOoIfu03w
hTDUoIrU6b1eR8Y8zoCzC33a7IEfW9ZnmUsS+9gs7vCitPvFXpWeEBgdOjmFMOYa
vyExtx12iowOr4U4GzmeAcp9LLl1vcF1NfShSXbOWAmYJI8Jw7PwlGG4jBZL+21b
OdGtePRq2sZMOhqBeSV1mF7zpcP3bJir+jI+KV7+pmYyl6OFh4zUUzKao5iGNuH3
5Kf4K+h3uYLvO7j05rsMPPIFVT2OXOggidpf3UpfDq4C67O8EIgV0KZdKJALFi2O
9icz3pEcp4gDkRv2qvXs5tJzKZsOerB+lY77NlmgWno2weid0nADWqC+8rrZpDe4
fwmFjVJCEyEYlnVtq9v2J02fN6DmTM00xKOZQ8ETyHWloH75mz3UgeMo+3/IkNO7
x8xexJVYStvgPpc9VZj8BvU1pfhwqd0E6CQb3tMcbJSaF1BfU7gPSY42NRun7kt3
Cui50OD4cCXMR72a8XmYcMQ8D4kd1d50EKaF3+Eq6I3YSMixAoo1x8pkVpJWiXgw
1R0XuJpSy3PAATOdBGSTrxGJE//NHnmci0/gHT0jlCI+7ABqQT3f4+7EyXqiUkiI
SMzKfKjctUw+q12on52o8U3mlyIck+Wn8TX/VjQSEZ9sNONIITd/SzXW1i8Woy65
l06rXOie21xOZGurnR/BZAlgvl3DWqOLXLpqtF3qa6cOfiRlaEL8MNOjUu7QvDH2
NBeyH0wmRnSqL9VaHnPZRhpsU1n1yIG6RidMfBalZGqNhPUIQqXMOYd950O+y3k7
4YUZSIjf+RY0rfQHMRsMF/2Any9OFMWBqykjU6mYEWuH4G9sIAfLj9JeGkblYmvV
bSwKNus28j3xPYjeO/1Js3Pea0OKMW0ugGjLtnPn8gtlMaMPYeSPW58fBC3Q1kfX
4xoLDaFBgTY6GCGBesSC5Iv/fQm/3CYXFDWXQcExDGt0DqCZ8BH1gw3y4eCoQavF
k8b1c3jjFdwDFK6oL47ZuArefciRKpX67z2sHFWq22FTUFJGpUEVdCvCLxRKD/dB
6EXkOCNji9vhtw+HjYm4IDjamJTpqK8D+qCdViKD11OPtZvbrQYvSQvW+Meka9W1
HSDGaA4fEDkJ4hXpJyGdmcH0WErda7GnSm3gV5UdEh2nd7Kgbs9QZq9GtTazQnkS
fiwAl8D4CNnTIlQJE+ohgb1hLwSrFFRbvDguG1idTma9zEbaJvkP5GbTUoLxht+a
AcfTBZajkZkm0aEhch7RFhDCu9xzaDxKCls2GvyteSf/aiDI3okJ4fzfmLyqhH0o
EQ4MDMlH7PjeTGkLktKw7uw5CJ4dBeSr9Oz6b+5wDP6sRYRtGvkZmtfN7eHkwU60
vt4Yw7P7DuidN754mnwld63eWb/44gQmWdLUSuAkULqbKEgIbvdsd9AtgvNnR8Li
YKZUE7zpGmkotoegmXw5ZMMSBWcjatvzDc+/45cHYuDJTCZmLPemwga7PlMhkmGV
HKuQmogjts5h/ZHZOHkK8rkj1gAihh9zdJ1b14Rv1TSaWnykVUknfnio0c1oozt2
9Oh/eyxDEBenlpy/YdNhJBjr5rECQiItvX9fE1gMhkzEoPzQ8fUf94JCbh+VfEBt
9k+Vt1w4+SNNO5i4HXOGDlk53GPNo/ZXtFJoatsy6tW/mBDWPMhjUwKd3P9AeSjj
6ZfRE5t0UyTmLtbegsQrlTo3slrKkiGRE4kXyPSMs+fBL/IDc0B5HTvKRBaxIsAm
0SPTkCtuVVZAp3pKcy41HiJo1QyPmtqrdgEPJ8jjSd7tglwgV8No0N8ofhi5igwp
HAGtBc7dgJWUKnutyYl+w0IwGMXUNZv8Lw8nuAXwhLCKlVFPbtsovSgAqNpn72fe
Q3Z7eFFfEjm8zF69yujfzwOHCCa2o/PK/pezRdvo8posxwXKbTr31CLJQ0fMCExk
Uqnj8CWLcWbQcLxHTI75vDYLdorOo+kNCy0ebh072F9UpE0O2v/Kp9KZAolCLwJk
5BcflNZUPIl9erPKEbwrou2oIrTeq/fEQRhMW2cf2deFFoBHMfcDlglRXS4QAauW
08gRDTJnYPAC36kOhVMYaKccow6EG3uK9/J+9EOYV6AIgpUZWsBNGE8qRPiPM2Nm
9JMEm5rJ2xXTP645EaH0MmGNLhBaGqM5alc/TxGeneqG3WHLJH7vu1gIwVWO+PaZ
DCJKogNWCgv2KGUnCkIn3Z726JECpGTa2Z5SplMHPYkV60vJsSZMBygT6QRL25QK
K+Le7LQGakEwY13k6fQDJDSoFHk9ZIi12nYtwZ/TgBsdT5osRV6EqLjXYeiz4fyy
34c83VXum/o9r0KaiX3OVkueGu6UNVPT/L7haIyo25zxEqHZFA26C+3xAAx6KhYp
Sa3sglJJhc+DDicwIj7Ojn4R1ibyveQ8oP/c8vYUxZdGLm8AfUEQ3Nz2cMOSDeEP
A/H5Q34wb35PzNKZDuS6tzafH4IUJxsl5RVFkZf958UfxRFOMjtr17ckbn1Kj5lP
80YP+yT8ALJwi0xJ+qi7qipLZnjQg/WF8jXZ0UEUIAcvJ4+JNEmTsAKqpyT8cKdl
wpPlINgxg8U0KHMRQx9qcrH/GRzYLaY17aD85me4b6w0fXFCrg0FsnJuS90lQLV/
nm2qjGmG9l6CDqUIw3P1PKKjRIpFqkNHRGbEQsU3UAcYOHxe8vmFcQj8U/FBlkSj
khVE1XHH4WS7wxnJUzN1gmKaG0KkV2vS5y/SNqweZNRmPFLbjZLrNIL7atBIn/+s
q4WLw7AruBEAWNtolLmCsbCIzpWhVuQaAqEofLGV0kkwLlM/OnGJ3C/aDjL8RUhh
ez1JOZNzDdYdEMcei1p3fIhusVbGKzHVZHLNzomJPryuMx7cGZvEM2stnX/owRBL
9SfYj9IbMATaiWeH+nE0Q7FuozA5/m3oBLjtazewInH6ARV8fTJO4B+Z7RlC8lwa
c9LjXbwGvaBP1KL67CuGFrvPAVTRVxtV0YS5xWaCGyS12mJfsAdKNxs4djbGzKM6
/ZowylrCmm7t2DXI7z9fRqaLZu+FmKD8793NfG+tNp7XlVlr0DwXMv2W1vguG7ZD
FJNjPmvlRzNcJ1hpa9makqIXgAzzW/9PSPlpBhPJ0kUz93XcVrHc+ZBU81Lyqpv9
cVitlULAwpnwiy4M2FZKlv+orO/TGZCYxqGUEQ3j2NZweZKhByunb/iGSAUPLdgs
XVrNK3MYxC5pLnzPvQIElfITADIfyTPm64+823wiigFm7fZ7oR700E82c2z4leKd
8fkl7P35G6f4QeMNio/DsdnGtcrjsjHjNo+laSs5o7NrjlAziGl3p+91dWc3eBYF
1aojKFY7pJrG+n53/lXttyx8eJqy5rtrR033tBec34x+bqh6l+30ni/Qwk426OOF
EuRSHPuUz4vioUOnlRa4tBobCiE7zcdcFC4MGqD0Jwte2bIfxfRXYa9UCnoqKKRW
veDs57LMNQcvotw2WPZkaJS2YQz873oABZnAErF29KgH5ljgmM/kTNUibBo3RBm3
44ELojzlD/AvV9xUoLlpwU4Kr/y/8qVY5j3vwlkdYyO4nL0yc40s9FrVFKQt/Qjy
W2TgMRQvpu4Z4ndtI24skLGkMsj55v84ln8uHpcmGvryZe0Ee397DGzAz8/EMnhM
FUQVOOyQWkagvG70zWGmKax7zfT7d+bX9b2dH6Tm268OEfEGcrerfWJErgSz9auH
d7+eJWU2ABA+XPUsLX4/MCDjv2AbzXGzrs+GyOUnT+l6LtTFv0ZysWrA2w/P774J
q+quZ5UAcuNrrTDd7y5XhZTcr4xDjhCG/hBkj4r3lBEiYW0GH16FwcUb+hZobEwl
jZQifq/2DScMNClBTambO/T5Rh4YsWTDHXQ0dRkHuRZ0hhUAlbpRgZl5XBEV69gU
Xl5rY4RXG8C5QDRz+nph2G4UqrmUxsRjNefM03ELYb+Q0jagLIwxmnVBhDhYFGxV
FR8PZWZZ5YyzfpFhFjwFzSJJf7z2OI0kYoTL8caP2efNS3SbTO8PeBvnPxQh/Ukb
SVr/UMO/4gzh72R6FZKRxJC5Od1Eo9bA/DaTuutmXybMvmRwUsInC+0hlA/xoG8D
uCveYGvi7a5YH8Yjse1bCwIxXrxub2u0BafVxZ8rx1y+7VAomL/RwQiDDKOKdq/A
nzWGL08ZuVZPfpL+CBX5HiAermJOybnqpNQanc/ldTofsOgXcNa5ZeuXMvr6Thy1
lBpiEwLqZc1Dk1e7fvkRLxnPveVwWB8+yOcSGecq3T1pG1j7DOZEHbboG5UJUdho
pkWAEPdtMwOwrEP06u3JJtzyrutQFLvrVel3Rej+El4SJZ6QzYRI/wZTTUxhBdbB
JoJWuYstTRGZntKIT58bHJLpUsXAfkmuXhwLJLGEBX21jdVUh9y86UWVFrUipKiz
xLn7608e/UVyBTFjGBwNwF7eE7af4rEzCsOEMotFZwLFvqe8sewmGvxXrJpNCETN
BWLFVV6E3Bl3uYopnUXWmGIUS/y3scK9dBN/67cKw5a+AejTFIlagIvONRhCFDzU
IECcLXe01be0L6H1pN0kq2f8klExi1QPr/SvlvDz+telphM31wHKTVy8Nl6DXOYb
QyaXT5+5ZubQBxiIim5IkgAXfOzIzAkHYALwtiz22zH0F4QaVN1wWpPQixJteOKA
PshY7B6wtcxiAwBlXtQK2osXtNDaDlv21FgfTQwFv+jCaqfvu3K3l63yDvUI3s67
AmQkLwWq49hLwgytBvAumzhChS4fFFSseRsPVoEFP5ivkksRNOs3KrGjXalGNbEX
SVJHgaEcrnkvscdKVkAWyTwr77Km/dGFAEU+ztS/OVXe/9uy/ZV5uddy9p2qLnMT
S//S7NB5IAqNsidWDAMnSYo8dbbZnnIht/kechtgWboZEHoTdZ7Wm+2mS1rlRBpN
aooSRsp+fSXcRe/rB6UFcdD0Cci+5DoHZ7syqTHN+823/uUXa33fZIZjMGYS3iZk
HQ+PhbL4/GiY31zkZ0tDL4g4PxDWPblMuYvqUn0cSdU06q5I4yEK1cS/WMclefDE
zQ9BtfoN+sNfb1HoLL2goid0OPo8cppZlgreRF+1WWvMN+oM7Rwh5ppMtJ9XmuPV
RyLiX3esRh8VGPi0VtosrhvYsK+OsowDcj0W6nof5OdguCeoFZ6xkLGFFqLrLiv6
AT4NB4NtRAw6oXUn8GqWhp2SUfhR5/Ni+zhmTNcacys7t9Ao5y0IaIW5Pc2xGcaj
3nW8+A+hj5GkiyeqGj8ooxtbvrj9SmFCOskbHtVtfdFZ/dQYgX0y1TsyeULVJ+rP
jpd2mRqko0KZCCUJRkdMUjhAbPD4UThIGBYOkhrSbbmPCUgYRSWR14OB0x+m2pQs
nrRSqPL787f47zgGY3YfibyA9lAdC1+B4DyQmrC0P6u5PKV76xz0otnRr4POo6of
eia1cGyKJ7YIYnZAo071bJJZp2Z6em5HdJqvEY+Pv8z12BFdI/3wgRRo1xRhHhXv
27JJ+ARC+sBcCca3zWUtAnvIWGP5Fj9flIeiv82m6X+cCCKl2OrH8pK9i8HL/Fp6
0NNF4kdrzKdnLJ3izWB1l1Z4EtOtnraY1i1LfWNaJlVLjYbmLgMG7rhipM479I05
vPpD+AsnLgPasBcn+OW2bH/JHF0qvZKQ6+U/tHjv+vstRYv/9NBRpI65kKYi9RbH
Uj/ryZpsPfnNHOa3CLhfCumCetF878wN3hGoqC3BKQDjOIr//CwDLIpfPZKo+Lph
7BiOwnZtdLGjv6bBtA6xRJaBfivvGNLymn+drPVKxHy0XObg43WjxidYLnLPtHAa
55AOEhx+rBLEAETYVXkyKBghuqyrYn1coom4vxVWPs7204nOqJQK1zgiZTL9Puf5
82JOH6xAAnp+HH0MHwznvnNVxTqnBJVf5r1UYyGC5JG7z1C2z4HPWdGgKKaJVzfh
E2/AUbdp7ryBWeAHWvz5Ey7MA5Le/37akesosZZ6hyPI4jdZF4rmutgtA961VRX2
MJsMpbds/z9OBsPsNwNM62XZyV22cEwNe6Cjp7ylGdWACArpjcLIx1pnGxeOajy6
+1X9qn1VNJ8xnw9O4JULWZRwfSQQ+hNSRPZgnwKsO7GwE67wwy+q2+dXNsBeWwS8
oKGgz5yf+u3wTdYexKcAPsrEByYKWTqZNvqoxGjuJMElAa8WzttZr3OxwmozpIu+
SFBnQCRy/S+n7CdGAVyeZLSsDHf1ajeQhq2ijFk35S1ochbwyt9b5/bTtF9rqxZq
m1yAwKW5o31atcnbpv8HnuU01WuvI7YXT6VIZAHk9J2AnbJSgqKmE43/qg7kWUN5
ql9teW4UnzinHqOx1UX7oC7TLnSnmqyEQtpTsHRe3/T385A7bPsjU7Pp45Ge52KK
yUS1kJw0XYqGpz0D/qLJlfusOIOsuet5bKM8ZK5QQfjATCZijFnjvU+WL+Aw6Ufo
tsd4krxSVps3PUnl75W3Kks/54VUri2hH/2PGehRM2xv0ef3fjbKN4Ac2IYbVNcc
Z5IAh5Xg8lOVF7MgoAQyqSZlsCYo1lAVt/yrNb7clygMtuBzJUrncUwf1fNLFEFo
aIXfbf99o7zolGNoZ9REGNVBV3i00Cr9+qW82e8z/pQls9bfNinIkY3jIq6aJGwa
QJ7KY9hg/szzZo3IcNvhnyACDlTr9Vs05RuYvaMBfF+nD7tbVQsO9wF2AQ0PEsPR
Scn/NPlu6bB+VkYo1YUf1x4UFc/hhyYM5v9IYmcWVxHHZmT2/bviiFyGZbnugjUi
nWrRB8uOgp1ADfq3cyNVuWRAExGJl3m/JCpq+qhQpexSKghqGjAhfus+4CH47GKD
18I7ABcNiU4WECBccQVIEk5VZeIjA5a5wc5bPoa3KmhwEO2Sna/QHAHFthWgAcsD
agC7Sff3qK1xO31+ejmvV3Rsyf0IEJ+sf9kIz0pw877EH1NPG2IBG4T/nEXzy6Zh
0qErFYYBWupCmwK7CMpFirnXLcSCX/uMjYcYGuo8L01UfxGyfbaDAekrI4NfXR6v
hO3yMvWNAlViXw6jXVYeXprcVoVaj3Fj4qiiwbzZdIn496RDUBveMAQ1eQ5mffua
a1wOLi24H04N0LAX1+2y8DYeB9TMqHFM5qBE9rEEAA6E9PaHdMAnS3zBp00mV9F+
/PbYY0+EYfoHu7izvPyEa7wwBSeYcyWqb0FV7OD2Xas1/6QBG6OZcx6l/rf1VuX5
SnVVj6IIJUFvehgy0idCsDsHaIvJhXQLXHRGNxl3KM4oKARTe1bmIWqyY1ynTMW9
yjXPX5AV/2ZVf/pDz64Q25RkBBJdFImDv7//NXX6wV19b0KxfFw9hh9csdNbBsMu
OGtOMPqaNTKzJPAu3El2yCr6v53kik8XEJKiUuroM77e7FHgyKiICxJNJtWSoJNb
ID6hljELDHSnXGvn9B7KmaPXDXVO/yMeXMLGHpK5Qar/qC/eS+EmxWrWGKBA+wIU
gNXkGyeOuVSzVBjhUBSvkU9JmPqD2hmYZ7ie3Vupf8sD7EagFqCOr4GNRjN4uQzR
8dtCyHEnnAOf+UcasKhIu/1V4q4Mq2w9IiJzo5O+iLzmBj9Kx+IH6qWc2Q5eOmyb
FPgmSmcD1KlllLHNMe5U/2O0DHfiZyipz6azvWLJoAsW2P5A1NXTz1Kd0LGXKnMC
09Gxo97/E7P4ExysoxVN77NPja3SKY/q3ovZV+0kb4ZrbESOcHsRKzJAya/uxVgm
oI3L5ELK8VsgzjQt2PqNoTDFsdX4to5rXDF3gYcD72njF8appf4Y0nrcEx0LYZW/
OiMTiiYJH9O3DWUICqZnS6+TykErk5tOUqzjPULNyHm3cW36fj3+VkrGql6HDOyA
SPwi5A3TNlz33gDrqEDQZJTl9myKCHSkMwouF606SAeJzKLybcVsKoFrmgOWdi2G
peHKydG3J5GV5+QdNnjR0i9OHVlWllM/os4uwNMjzIg8CuhrT1Oi8xSlw8cPjt12
Fg+sKDFhLH+m2XsIRgeWmNucQSfOHJRsnAADZCI4RUDw4J/JakIULMIAVgqbdTf5
8bTdDUfWC0mNK8bVld3iHRX/3o0q2GL8mID+YNuOPVjA7G8zdfNPCWPRkbMqBLu4
VLpPGqruNF4epJVh4ULCfD0cpeLvvFxVb4FTm7btdLU4Y5che0a7MavhU8M3U7C7
j/qWae9wi9BcQarb0+HETJYlDyJOPqGyE4BW+8YgmoxIXvxZu3fP5GSjW7JNXNJ1
GWX56JNd6lepRfXbPfZ8jHwRgj8bY9vI+ghjUvEZSJMPKG4psHdySfpGOFJK0qgo
iJJjAVCyyD55zEdsb9yx4vu77cvppxSB4D0ElwTDJbtXWoZg88Y7gqfEEy9DnJ4T
ztky8MJYfiMuhvpTKZsp2wReo21g52RnU88IMqxYqjDCNUzBHQDGeD1Zkdv5uYnB
jRQ/+r/A7bsTL7diN5fn04K9RS8CYVYd0r0BA/yPB2LczhcYpzAh8EtmbiuMnrmf
wFlsP1Vj0RTtUA7oXP+MTSsCF0fbsIK0FTJjkz9Xv8wFFPg4gQIid33kk1sN03yu
f1cNAw1LaLPSh8g38exfN54FP7QIUEcNZrBQdTtIfNIRgPMbHWH5ywp/I2+QBuxi
7RkaxHevLcCMjRvhNcaBL5Nu7gWk/p/yEknWImkzdXmXoxkG0mPxROtVd8+Umx/7
pT2ePc94y3vM+/OFFkKEdsLzaZFBxPtqUCP5GwKceU7wFAZ1Ap7WemsU8jdVDKf4
1fEC84H5KUy84gGoVEFI5ut7yJ8Dko3N646EwnJow1e/Q2ULNRU6AxjfW2LmVuUd
nW2f9ZKIY1IxoGAYkDVfcM+tQkumTOx6YuRKUL9zA2EM/vl6PZct77YczRmAdYNU
X98OmsdS+JzprMmaYWN/X0LXNlY57XT48eN3H04VMy3qv8EUrE403+gpC666wYn9
bkuE32t0w/iOloXrjhMo+08fAKTn4hW+cZqvpmrVUmIv+ulu5+zy/GYzi9x1jirW
FPSCGhsYBvwyGI94ckq3RQQgaf/XvkwODupXdrtkOpRE6BtKsxzzprYomgD4KePt
tuErB0ObYFWSFqgQxpvAqcPVquddtd1ojE1bMhEuWolej9t3T/a+b5REUb09ASIC
jqNbBm7UThEwVxqBlKBavQn6+OH0uNHu232DkH9P6SOWrg0lIWdl+S+Du5ksoHAd
/hqGlpoon3C21SwG//8mbjZ2D+KfY3epfHMLhOUG487UA6u7pkMZLTU8/vM56b6L
8pm7IiMDFLiqUIyxisg8cRi6B4wdzhHcqxeoWnUIF1TvOl0iqy7v/ucVoalPucBf
0g5Y3GOF1WSBHQe5U99d1pi+DXWByD1KTSBvlLsU0A0jNYdERrJaV83piwz9gMi2
sW4eOyiCWb+jokf823MybDJJ3SpPg46VmPXzqmRSf6YXffB5n3smjtt3S9rhmPR7
DdxgAitWHUwPMtwIRMMmNOSkAjeAZdc1jgapyKeF3em/jvmCGz9h7Hvhk+jjlz/z
3BllebaZIVZUGQ1nsdTW3iBgMtLUYLPhkjF6B9byfwDh7CqRdgIH5UeHq/DijX8G
4z3T9cMQviDV+gdS0xfpq519jsfuO/8kIrYL7jeWgzmRNXmS3z+G9Vo45wQLku1e
VTpRpJZmu0gdXscrTP40vtFT7n6UKwkvZHjhT12rLVYkEn1GEQNAg633iQyPyGgD
cwfAj1wtWQm7WKbGQeYvf/oxk8gWaQXBSknLwU0gG5y5XXsytaLSFiu58iBEa+9r
t1TZXHgdAmLekvZgBeoYnRA8n10W6fP/OTIpFn5aG60MP8dhG4971fZSnLouXndi
JIwNjSbJIxF2udwLiFvLHSI/Lkvb9FnCxd/bX8Dn4qGON5XHIsWDtxK6/Bh0yeWg
3pVtb8gXXmacdmH0hz4jJm/LQWocr+MKGRIOhQo4xOdk5U1QsJgjRXsnngL2FG7+
KQwXwCms7vNQRWt6G3rsX2uNRf2iCYhpkNbpljjSHL55VTV2UIXBRUdQwo0i0Ppu
SLBhLlAH7o+2c4C1q26Lq6hEZ1Rn32VCbDmbST7SF+UJNXm+NiCf0NPH8j43BkVY
71p0eyk/6tPf2o8KSGTwo0K5zh3CeUmkBkXL1XuNqVmaCR9W0fTAbZaNQNveUNPl
XXWSM6m88420DU1ElwA/+gg7bFDBarwbjV2AdzKYRLR+UN6/Ln+kYt+VyC0m4afh
RFxy375dkhfdHE0VI6YWueI808dX+1U05zqKo5kaO09jbHERGNy6zqHahGV0y5TV
cygfMst6EGMBqOkFk3zYLtXbry+T0Aav9grhHLmDDLz1O0ZiRMhJIbzpmnkcyQDd
wbElnQYRMY54/y9lTRmXBdANxJ9Ad4pSuAfIawh87vS7hZQ2ro7BC6rq5W6f0K1O
Jxl+T4lqDeZOP135FK5Rxu442GEKhLAOZBWe9HYVcDrBNq+Jt1LZvHodUBarIVCK
wAHfbXk7lJKI84FG8v/s5VKfHFIXTzA+pvITU8YSf/QJjSDmfoi1JM8y52FrOjf/
mI2HQJkmuWoS7caT4ith7g1pAyNZktLmnv89zy33hTWlexhbEV455036IK1I61gs
JCDxy0WAp5mGE+XZ8NfPyFa34U+F7tfJMOfcD+pKnkQod6NuhmUkznHZkyu8inEM
Wp6sK5g0CEZco1FM9Me5giiZiOt94fXqOWRs35preBWESg6Z+2F6O3+OCfFSA+OD
rpKDydObgUqBvfROleih2iM783z6SgfHD0NfBdi2wT4CYWFcnGiujhgxR+oHaLRc
h+RS0dNDwOgs6qeIVLUI62xeQVRKm36dv8/q5iAlAN/8I7Z7MkN1/QeQj3m3qcjf
Q5rWO0tWjAuGyUsVrdHLCmXMWMgTMt/LcV50yQbPqavGiwB2zIWUmVoMEn63HjVw
JieAUHeXYh5LEf+yiHcUE0DLeIaJ7n6shL7KGPkwAiCtkx+MsPU1BFDhIDEyKI3q
AkGnXNNoLdKERE2fYoo4Lb7gpVaCHTYmNsAZeAUTarXzyXB9GvRSDDSkV86bi+e+
blWCa44oZP+Qe7QUzGYRIKVz4YOG9RgmNzQJZi220sfmeYGayS5T+x88bie5xgWq
JSWi4AQVfoLPSrtUQP93SUjWogsAzjJE0XEf07SzDFJFfT3UgCwurT4LrHT43xaF
N/sbkW6y8/W3qYg2xe0lPnJtCGdUQqlyM4hZSlnBK0GPJjW037tlDP963T6bPiFV
ITHSo4b1b4ncC5Qx5GYRRsTj97LTZaFHQNaBpXc82VQzCehcPYGx5s9kTf2HCVo6
jLyIKKMILMkkQDZkjOxcf4CsGZqx5l0JhvbHqgrYhX88Vr+978jf9N+Pha3hWZ2C
6BSBEi49KemTPruSeUSAXmMrykozDCLu4y8XO01JKxoM4AeXXoEPAe1MFUNhege6
zwhGdpjl08Pm2C4Rhl8V8YvkLBQwFozJlCI1GMEJM7foSg5W9y+WPUxLygpZdJQ/
uyMVZfajamSiihSDyriLyOgJQvU4xlnzpOaiRfhpt2TOjaBhKn25oykFZ1kZ0vo5
OQLGEI9wbgvDht4ZasOukEzACnsZ/DEMWSEXo9/6wGSndTWb7CrEsdDvcZWJgcQA
xuW3cECCep5DjDArWPoLLZGNf9JLwm5GlRFNUGTwqPaPKPhEQMPNZ36z4sQvh7PN
jjheA4UG+NhApbpmWmnlsCJjoD+ov12SRBowfj69QbPxR9Z9TK0IJ0Dr9Bz6wzdH
SaUk80t/kkbY/J0VLub265g2NLjojWqUTAmdGAwjeuI8ZaQI4OHfNLj/CYQDEV21
fgVgdf+PPEkofGbdYbyhhosRygatxRMDW5T6URRDPS8nZakDD12vIDlAfmrP2ibZ
i7b3xLBVjiFTrpom4cm7GdE6N9W+uunqg/JOumtBapLfI8GsFO/UqdvFqanFcx92
Cg67CDqWaH25Uuk5YhUAHoZN8p+hwsblXmstndTy16A4qOEqNudNQlYGtJjy+kpo
gkQt2WlRm7bh1OzmkR5nYIWXwvCtRuYNZ2u7C1BhJo1Tz5dl9PUFgX/tzB4VPS2q
N+HoJ00111WNvpRbVbz7csQiwKcLeZohe1PQQFafKAYcyNjvuO054o5RP5VcvR6G
A+NOLefIr46XNaPRmfQIGKLjhuKlxeLXO7DDNxACx0Y7Mds0xu4G+//WXxPXmcPG
6Ow19d062IsX6pM7izZAdSh81MScuSf/PU+ylb7ESbIEhsRwtoX0AjUQIusQbQ7i
bE8BBKEQfbspzDEkzZ0doHCSmgKhFWUqIlCCWvwy9bQTHBJ5yu8y19PzML9hTh6a
6cbpWnCaDDr9xSco8GGoqApDlAv4er5Eci4V+v1083IzTxjaVPxpo0PL8XUk7jCt
y4xO1AodGyXifqGM3NWMyZpTeiNp7S6HzpJ526fhYk9u6OP/H4iqZ7lbVOYZysTP
b+zR8+owhskN5II/MoyTLshtR9AJlpzVfv0eCzpxo3ooWrOTTd9LpUlwTv/zcuhO
ebM3nmDeuzojRb0a4/rIMZbm5wke30CCFEsgdj2PGliMYWVq5ue9TX6YhtVkYdiT
V9tab3jUJrJaQ/oC2XcHwnvBFD5iQJw5acnqPufffom78qqKXVYvMMBVuOCXKN4g
bxReWM53KP4lpKf+Fez02fIJuBjzuW8TP8UVq/mSygc/OHYGeTBwhXu0ua+DCXkt
yI5tDOJ2xjPZseBxZZPs7mGbHO47MTkvhbJTHg7Q0vUdxN3jqoK3T3ekNqbItdvw
R6xmlIH8qRSQKfWP/2dAV6f4g1Vu4loZpwsf+N6QaMmQjx4LkMQY2duh30T6iEal
iK91WAg0yw6dushag8bd5csvKE+4wJkoEuPkaTRXj5E7N7qwPIjQ0UaLq5/fJeS5
viWNqeGvLy8c+8WoLUk/FwmVob3MnbqBTDR9MUnS1c1cvoktKLkd9iUYgNNedn06
63I57nYoE0ZvL5Vt/8GKJmMl1niiHsoTl2MkhVvuiqHcKP0H3rq/fhz9930gxlf+
sN6IsajTdZh5zi+8/SVFSB3dX4Iri5qllLQ5+gx8ap7xFJDo2czYVGTZiuGLkUcU
c+A2Ut2MXkj5xSTMu0mDArCIN+cou+dCqYJGJyYTY3UNvFOTgmcF/KVIKkGoEVdm
ISyvuErBjrasAvY7cfDwhJpek2hAfCkMePg1hkmiGFLw1bfDQbDlOxDzqjlBsIVP
dQlWGc55tevMoE3uKOw8DzjHf2HbbGAmjVGlgkUduD3637uxeMURbQkjFS8xW7dR
ZfHUiAV/7D5XIa6H2OR134RtaR9y2+HfawzH1iaoapeHCQM1Nsv7LYTRsT2k2L5j
H4uyWwXByhIt3vYub9lalVZsytrtfK3wYSYg0b2s9wo31VsGv6lA9IHK8mrLjZgR
0gN26cgqmAJSnX5sNzEnSVyEzCu7SEVOD0W6OuW5jEOwU03kKAhPeUzIq+Q/8Xff
kUzzms899yzGGb1MvFOy235PiHvOEiK7xO49FlPMlb+XFqa6s8H/mDe86YdhC8SU
uhwQ+eYXON6kBgy02aj7aR0liHhWBJtvYw+l8VsyBjCsDfhTBJzvryCxqSc083qv
PIwgaIQRIKPbw0NweWpklo+a8IMlVVkTQCfYhgE91cSuL3Cq4KQkyhwKna77UVS+
ZXYa43hGrUS/tSb/9QF0EWF9vfoskTEcerVqIu+td+EvNciF9gdtD7uwVIzHjt3V
voApKJOjyr1bWbUOx/E0bmdi8JFWFnaOAOJuyapdU1B+PqQj0CNtHrmL3OhTfJU1
eOboCTmT0DhJLhH/HxlnWC3DX9SWIuYYrApQzPrcW1RtOKwQqfQSqXncFu2PKT/S
q2MxBuVNPs9aJUsLdzvFz4+vfl6+q8ZqeyOy0eh979YwMNNCVhvaLlRsaSMny6+i
yxDWBBk1p9/xDSGL+m2RxB/Lhg5hIW9caS62iRpoLIYYwIUB+Jd5UU67lNigWY7t
1HaB+seke4z9ImsXIkRLmS9/wUzaMJKQfDqHCN2Kd3/IfnQT7q/7Dfer63wxEk2u
OH44zznDXKwbwV2ydx+uyqa1QsdrmcGUmEN+9sfBp7kQqPRGS4GsCQ7YGnb8T54u
cGfe6Lqv65vfMH87yq0uqriHlffZYmJjuR5vaNqdbDYRsnFiHimIYmKcmnXq+Ihs
kOwUrLCReyoZrYLMD1lls0dQt7mlWAA3y2Ye0ykPZBrNwsk45nVOQBAywKksPO/X
mpAbEs2e85NyeQliOBaCc5l0vjMEszvzktetp22JbOuMJrE3lA762otdwPL6SvXC
+yRWTbygHZw/2JsKboCf1WCjxP4FeWeXWRA+MEdNkqXeh/UPKGIRDLoUUA24V3o7
lHX6IsI0dbqUa0ly+JxhBkRym8nRUmeZ+I9lEFD5DVACLPHeROZQ8eV15CDsIkC6
mJ6e2bl31+Nzt0Eb9ePUEinOrH0e6tVBTiz8jez1P4rIEliB2muhUwmdwaRFFwCY
qANwZfQ653fCn+s5VVRzH8S5r4V6CUwJLq+ysrJLwVdJRc4thSEzQsRoPKe9NGKy
1jiZy8lJ/wWW4XreHmiYXB3DuACthHzP+l35hBLK7BS301Y3FR8hiG2pnXSUrWDq
6YFuIbpWRLDnmoZuqblDVy7QOqtmFFad2Gzu963FjPRsBFnlpN7U3VnlPLdz/TB8
p1r4P+Vq5Ezf1y/l+LUlQ55N3ryiUeOk2vDLLUPyeFfwhoz0Z7qGuy4W4kGbTrIX
EQ8LEcIdTK3H2ah5ad4R9BAGmAuFbm+gJdwWFMjGQxaI5giwTti1q8kDVtTR8vB8
g4N+ZnlAfHiHih5Phctr3xf1IDFS0/t1pOkDM8AEdFp/VLO21qXxEAHePK8PRxfb
M6Tn7HMw4cNdAvmmJrzrpExgsvEs3xn3lQafjzSeuZebhzYYLBXMuNr0DsPJvmLK
tyxpIp+xKTkckkNRnNOak3oh5mC8K03bP4Dx6Vjtz07YOX9ziLQFCQrdIuboyTcU
CBsVvThZeK2Af5rrlW8PLvYI3gFYO94Loia4wlzWepMmmDuT2/S0PXTYLT1+2zhi
PfNUw2t3n5N4nY1c9vuDuJSPdmbjynIm0ZUU52jOWvvyu4d6rI2P5s3Nrk+hVQCM
I/6GDf7yVfjfPqMonfX/1NnIIm95nRAoDDkX7F9JNNLsGD9M/P9fZxt6bqHlunid
b5PCsJi7uAGyvdE7oJhfFn355cFe1Rz0ae5uhrBt0NlaLWDmnloBqbenYtUH6xXK
mZliGw/+ARnmHIeA6PsPo62mghoLMBLu7BLkyHZ60O8+Gb19lAPVCsq50KnMqp+O
nO8xZO7mo2EqvjMEikKlCdk3h4ZyoHQCwNFFsuHpxoSLeiJ4IhUmZHQHVVyP1V7s
PQT4qyLqIXa1S4IfHPxpXNKuTjyo5D/pWnTK9XrcROkYwRTHVY6rt3kUlEyvKJc1
C5bF9Ftclt0Kc04sFeOJX2kh2UqRNIBxPiw5wfd43JPAzQej2EncPd+twloH2F9L
X0nb+xYv8IHCiqD+n/4SNnIzAAY3Ocn1fVasO4J3/9M9GfFymi5GHipgxEHlbf/f
7wMaXBOmtC7Sj+BTgrIEXZCDqs4axYPZUwk166cupNubsGPkqmyX4TXEIahgiKp4
1pA1hjPEfXAzOcZJsLg97Q8nMUmq2rqimaFIGBuIx9BhJeMuPWDbGZ07ZBalW+4n
UcSKG9TaTM2OsZhXBSYpefXDIriIxe1gGLLVlYQtO+a5OxeGDDk67vy9nXnxt6q3
thsMhAUJ8SL7q01o+YNizPphBwJg05DOW7CQUWKovv6hZWsCI3bPmVap1j2bXJ57
DxONwnmGmV9nbfVp9NBNs12+5JHpc15ws+jrUuWugtNwKgy3idVhzr1kgzFn399W
7NbvRjE4WlWdWYWVv8ZWm20Qk6IAtaSrq5F4+V98PBNMz61/Jorb+t8MIucxdqH0
qv9Ui82tZz2zJadElnvMURQhi+qBt4vVy7KjJOJ6lvOlGsD72Qg8lELCT1GWu3kL
jra455xXveisdH6l1Fp9LYO+pkvCHvLXr+u9WcOTIn4+9bBAEXinYlnWrS9perXl
r9GMf/30sFALyAA2zH1dvOvnWUmYKpfRFMQH1e/fa9v7VTaLzrtd/oqXdpg7ipt7
aoZ7eDCIg62m35MaC1SPKssKVvj125PailxzZF2pK+hyH/kfVkihUfvAHdEsX0xU
5aDP8GLdBPGEZ6hWxxfg1Mf9wCBHSSIHxenrxpLGPsTVBTtpGfefFYgC/X5+XmaW
N/NQ1u1dV1u7ehp0H5vNap0jeoKiCWo/LYy5hmsj5CikVOcFgxA6uvYjpNwnaWbb
tk2lNc6NXl6Pe+AwgiIrmepXspQ1rkg94vI0CMXQ7Jma1YsW0NRffJ/VZTrlQGeR
+xyJtA5bi3RhsdWVRDpwd1biAdrt+wLmBwkzTAreVF08lItA3rfFJBhYw/bXOd5C
IBpI4+0V4qr04TTKWmAYQ1XXtuqBM+OQ2XG1UTNo/zRlUkFu8LfYUEhqtxCZzBbw
KtfsTbLXFr5hUtNvJpVK4ItzV7wg/oY7U+LVod8gYFStzkw99ZtX3541wa5DjhNL
kQhL4ecyg0DiaD8db4rF7/pjn2FU4pEJRfvFeUbWm44UVavjhj57yK4+WlMJiHLp
yg/h5Nq1JKWzfXhKoQLgkRDPzv0J7ymxYK/QVK2nSMCDeG7MN6sUwFQV/IiW2NDR
mqOf/0Pfb6Z+1bm71G8DzvXqbnf6CSDzmX0IKUQx7d93XujfQBuvgwG5o+UaWs9C
7eYVgHa1FkiCTMchTGNxGewCS5ZPpEABTW0ojh5Rqx5JVya4naXZ9p+qy8L5326R
5ELRz1BBW11+QJ4NwQmgtePOZ7Cih26xTkyJMJP6h3TU5HfeiKLFV8shBuz34UVm
CH29Oi28qE5KShYSd5lKKalrr9qLO77a3cXT89hDabtG9+XnrUjY3VH5W4amIe/9
1tYIef73WiZ4s/5oGB3TOVWLNDWBnzB9mqyxco7yXT5rYrGpN3TMi4lKJcM+pUYL
2Q+QgJtgi5svHM6CfZdl/jClnGibRmFpi/RRjWVOPtGfshwHU1k3cX/wQKT56bVg
dDtilol2aICGUiUOn0IWbWEII21bH39D9q0VKkocI6X7dfjhO4taVUVvwBCpKZ+G
vWS3XaQL65TymGdqcZX22e+z12u8eIHbJqm3JSsiTNyht/TJiY35LFyJLBwQEp0Z
ZqGRdJPhUFY+uZvcNfkNRZHPnpDcFYihQBuIM1gpLoZyur5dT/TANC/v6dzuzGLk
XwNwFGjNj095bDS5zYUzUTLJ+yhZwAqk/ikHl29CC6hwRSwfVp9Z7lt2YVimE/3J
1g4D/TmGVAh+oAd/MaLptgHl3PQ0StQcmttEB606Ak1UAkjknJbBLuQLNtqKS6xq
31fPrYdLFxRORO/LdrwXk3w+Q9PvpVEPLkonKayd8QTtPpFdYBurpMie27CkTWsc
4uLKpLl3oywOOZVBfYJ3d5ZMBq/PI4OcqDLySkXiT9i8z8QQBQ75mUCyx8bwDNte
0femjgRy9CPFwkeVGLpNO9Wofdi9M2WzyWrqy0pUlRy8uUQg5XIg9zTz+v7tskQA
eBV/Q6l/xRDLDTr1FNESJni9KOv9rd7n8RZGd7vNCP89gb21eWRN6++NKlRzkS8l
onWnbIe20eHiHnZbVL68nex1D1OL0V7nT4go04TDn1g0FTvHzoEeLLkFlsckE/Lm
t5pzXh+fZU2JyXjFa1593J/kfsy+CQ14bQEI96n6xox8Udb/oGcBfF0p/KCEGfNt
rinNWybwJpCUlrf3/0VIMHXpgr23TY1W7cBIhoxyXU54D+g/oeNOR1Y8RdmXc5/6
Rk5qmCC5CB1Ol0cWbZRneu/ggxujKck9dxZAgVFaZJmhGkxS2w3BIwcCoREa7ikm
+YsezJAqgJ+iGsjpgZIrZw7gFUiLBuSbXmB4R8Q3+CrnrCA7Da00Qra66CL1Evtr
7WXq6hFepyX9ABwWaZTNH5cOsMPYeGJ7OYfK7BBzx6PbWXMoH44miqrQ/s5fcCsH
ualKO4Ci0gRVCFN+/6rS6V3O4tIslTOoX2ZdB/+x2ShpZZQf6rdsET4ClCYv+Sh5
ywxPSOBovfE77e8jVpXWy03NZMZj/wocY7VsxDFl8BxWK6BQ39bQOZ0ADh6XQHQq
R8wZOWQiLEJrOeAJ4H3+MUzzP5LXEnFvcSYonlesRxstGjaq+iJLk3hWCxduVc6b
0m6cfsswvq6rwnPTwaEHn0WVNlm43+BH0QRF4OsXh+YcP1WZRNIf1v4LbVB/uaah
dvp4w/wrokCkUNNrGnv/ZnbVgBIcdCXamliZCE+UxW8esZty+koIZRc7z+e7UYzQ
OY/VVBJ7fFBWzx5DWiccRukWL+Se2O411mFnyyRrWL5CKe6qzY9kt5goa4EybcZ6
jGx6vlij11kmWh9Pw16zO659tQj+WpMAYGNdG4AyShhbo8upEnlA4iJxgr8JvhwR
lLfFEsnGYmGzx8XhspwH4r82987wTiCGfHWMpv0D5HXrMdX8elWHSMpiz4k4rUx9
iaQe3KKF5etC/rxjWGurNZv5pqjdqpwqW+eMK8D8c4Wh+zV6ur0rLzbX34j/ACap
eR4jFGU7zd+jZref1FXFE6uqzcKc73DD7SRoKAWlmqdy1CZvOJEtm12HaUI8qs5W
YbnNTaidWY+EcpshfzkT4adAxEDV15EIRHL1xzSqBMsYdgYytXUYiLIYrZZDMaFA
yz6OaGd55HwEkx0ui+Yv7uNqsFXrZCxviNDkpgfuYQkk5JjsMe4zdA49FhrVMS5V
hP10SF1xH7TrWpP+XYYYkNzeHCdTvvksDh0ZkpV1lXDoTsQ0Y1cVm/HbpE7Xsum3
u35O6btj3W8gBu0ycgsrNZo14xYMJJADBzX2995A/uUaIqyzPbkEpDbLlM4p2yXo
dfac3hoaZu878PJ4cRdl0wcyov8xdlh04MhfC151WhHQj6uaQW023NHRbNVhwHty
GnkLXrKHdUv2ooc9eMY2qCzFbf46asM8NLMPcUUCZMTAMTHOboTp2FGvveo0Tv8U
XbGouNc6w4Tt5+YivfIXAHdNCMJVauPiD1SS9FEibKvfXGOl9vHBXWpo5qcsG8vH
8K4vLT6s0hr+49cCcfjS3gcOdYwiQn8siSqY4TuGcbPxhEXFj4r7sKI8rHptuf1u
qrJkWrPxXiWmAUbuu6qpf89BcrvnV5Qmg2rjocR7hc8caUtRXu/9KsFY4l9ALe6M
1qtkDMTKBzFYwFLEhApk4kxSsYs+sKLtfIk9pWniltfG7PO71Xf2mtWVHaot0V+6
0D2wdlSue7Y3vyJlGcOxLY+e+NgGAiGTel5x9ug+UzdyT3FkY4emnSKnHq5Fx/pv
53SDkk9V8att2gQGyMH1OZMN9n64yB4EVFzb89uy9WlkoRoFoDGoeu48LzaDhGb1
hwMUzIvUtYZ8jWHbMYNGmfBQb494idzYcmP5Ev7nG8OmNqOfRii54B1mQ4tL0SzU
5bcm2ZyNagESu+HxcOb8AqMd8ypJm5SRAnEss0Pnup2RRnEBRuQmAd5EkzvRmVjJ
wIUiuY/K/8LHCUqw4dm0FseAW0yx3S5xclYf+xDr0ZmV79sHETjJOhurFTfnUmA5
LKiCsn1rDRAeIDTCkZ1MeSnMmLJMj2eMblMBewKIPbz64ewPtAq9inBJHbnbcEOt
xSo9keF3g9uDU91fbLRD3axO2AfpRM1+Pr5mBFLJFmXwwLKtydoKHKC2omkr1gVP
E7bEIPPjPGA4QfVhufc5QYC0cgS4YKYYxxOMSj9BMCc/5SovjAOjiWAZanO97PdA
LAJs884oF27Spk4T2ONXs1LCsOhUrwyqXpMHN/iqr74dlfr5WQbOj3LF6X2UPTPI
zofluMcAB+gQxXQKJvyCicC9Vkmf8gTCD9FVQn6wHK1cBL+hXmc60yY+dxAE0Dfv
HHmuFXg+EtLYoSHoAVQHpI0utxZ8EO/SfOdJ02ZXObtDXDAfS2Yds9z1YOkKQAO6
t31SVb6Oyr30DN4cRVzBCYhZQjP2SfUccPFFxsTDzk5X57zqpOPjBp91lm2EUXY7
MzDvdQledrUI91cIO3uzajmJftBcZ6TsSjCuosbbv5fCbeoIj+nn9pzfJ4H28mQ5
CF7cXXYx9RINF9lTgd2dE8LU4anWBPDixRv6z/Q+DF9r3M7mX7mWDkDjvJsTv73l
7TQ9fkjJJ1wpGTZ7Qnnrupa1fG3a0Bmj/vhHGxcDphBE0HlFz9I7Gc4Cj9dz44S4
lkU8+XiuQQiO4YtgsJKuvT8R58nJ/X/UVV229vA4iDXfx+T97MrOAvbyA2B8yvo/
m/PYtAo37n4S1LJcqtGt8nWaVSgnUY3Epfo5TThSapvUmU1hNOWb6l6pyMiLGleS
cwqcZACAY8iA6rM2tQXXNBr7n7bvSu2yDyK895K/RS/oNEQHHuN++a6xtEr9MI3p
ajo/S8SwrLZlgN9XTxnBqNZgPFixO1CJ1dFOYoMcd0dUFLX1dx6RSFQbE2NzwVhv
zBa2Mt8RIfkq2BmqEEzxuBVW5ev+f85dmSma8BI5nrdQy2IHagGbI/5Mq4YKXs4Q
oUYPgCzDv4D4trks8fJagLiQdsgzkYpa7ZLx8O5L086Q8KC5SJ/pQmdGHS3YqNJI
B331Bb2WYZAz8ms1o64egEa7YO4H+Ohfe/ELbPmaP6DPZ6X6KWpLR36LLE6HqYYl
/UA9zHxHiUf9hPlFJSSHSpynlcHHX6QkP5P8JUo4jSzFZmKLqDi5n9x7fkNgvdKw
WDLl5XgQflFhk6+k2seoiCc/wETgLZGA+W6/q3XeyOh2M58Wkr09moazrlTlVB9P
kYToHrJq/yJmZ116HYcH2PX/SUOZiS+rmaIL1CRk/PgwyxJIn48Al+FUQwwUD5y+
OCGNwraIJjT755mOUdGYJSu6Yixq0JHKfumx8xPlm+GFlcjUX7kyzcokETjug4/j
9zl3jh6SBIWPfYEJcQR3JGksS4DRppctxMknjqsivpSCfYgj2EUyLpgaaZFcpdk4
PtMis5PBLv2EcSXsRnHfHll5jWToYkYp9nlcidYH/3eVH36v8cN+8Bse+pvTr5yq
kJkHU/JLdBJ1co47MkZWoYiVIqc9NhopE5lev8JryqS6PVti8T7fO+3KJUi8SCXQ
unQR7uosRpHOFbp7oECbh07ibjeFDv+JpsVGchFgDIX3wSi5XBY4dJ5aStuvzaFv
Fl6aLLw218kE7/XHG+1N/EaAC7ohUash9+EhRAT2sJdfunBA5evxjpA5zfQRgDLT
Raqgg9CxkchjQtE2Lnd4rATJAmIDCs6r/AXXmCRks1pVplgVvu+0bL/xujXxyr4K
FsAl90g4ApljYdTE8ki53oLXJkLZJkV/IauRl8UrBPEpnFAl175e+4tltV1lBulC
p906TLQT2Jyh8RhdVV81XAUUpuAMwPqRut7Mccdy1jp1lMttZ3eMqfbRpqTRR38c
BGUVJZtixRvFzlT83r20HPH4doKbcEV7tXf9T8k4yEBpiP7boG0zLDNd1wdk5d74
QwYULFU7qookw9h8K5RSQzME9tdqi7pP/2LPEKDyP2mZ0W3rHaUcuLleMGWWk0Pp
6r2W5txSzM6wAX38ag+GlW4U5RrPYYnph8hg1J+eJ3OPa1B1bZ5TslHjdvwyRHPK
HsdOWtxDGcPL+OwuJKJMwG3dG0lHqXvWmEKJ+oV3mj9HsG38FilQ/QjTknKsV+QR
kG1aUZH5jmXjR6YY13YjzPkhnwoG+pWb5brOl/J2wfRulgOImyZXf3f4zfVSK/o/
1iGe71Xt+TpbVLz3WSduF70I4FJEv6PsLk+GSTUSXTk3V6ekBNUGSPawj5e1EA3z
8bttWzZDd4RmIxSMQDrY+6QaGdXe4EsfKWCQpEI9M/DBn7Pk+UwWyL12GjaXAruM
sZu28Fnl2U6Tdo9rFFbqg0Iy6RbgPZ+0ZlUCZqxcZYakH8letNwsT+YsHYVksS+M
XkME7b7yL8+EZutqzt3NqNag5PH1D33lmfnStpFoNU8Z0VctV9P7RAJceGhNgcZr
IqQ20NfOPf/EVr9c49CE2Xk3Kf/EvXSrT7B52I/QR7e6bEoYUbcUZSLya+MEwHZZ
vSVxaW9mJK5DnJngUa2HH7ee3R1fT7WCyDqBLKKXz6tU+LTG1Pw5zQ+J0Drc1b3t
E+43rl+2GvrUjCDlTK1Acp/82ik75M3FRguUADM3k9AqUarxGcNOQbmctQADlXXC
pV9RzaL4YYaRa5STnTitxU+uE7CA9A4AiK8r6tnrpQXIqFELvlDQq5ADx0RPeUjO
YjukMQmI5iwR2EWlxVoFq0baDambGaMRN4q7SurxoKj4W2tXSmk2nVgM5pt5i1xk
Za4B3STWTwBcxzx8XmVdPfffyGnCArTQWULwexe9SA6Aps+IpkYOItsrQWK3VghH
xJg/ULVwWzo95IEPUz9m4G5+20Nan24ASyGwpnd4AyJj2c4i95xFbaA+UdGFhtXD
PrkAJrsTjnporTBysdv643C6bMTc9UZ9x9LwxCnBV5Voj2LVB25u5ct4KGVAzutB
lzuqYxVh0djpssPUJ/ZHkLnGwhrHyAyOB/gnwpEEi7vNNLOsLu8rk75lF40TluiE
WZGNp5qPIQsxCIjldLjXjC7T9C+2eQHAJydYjwYhK56niorEU3eLnzBvloZQHRm3
dsy8NYe2CE8ouFbaKQVg4oAxdg2Dueaxbyte6UEFuf3Rf5ol3yLAM4zaE6bOkPxH
dUHlWPXzLQjf1sUHsyKZrO8CCV1mjDJk+DZKe8g/5eo3WWOK6XfkH5usOJeR1CD/
S0GflicNm8TNX82iGdHLPJJLBXyA7czWrqIaXA/mSnB7n978dKlfqGOOtWYcnpOc
gIF7D1sMU/wDT8f5rsJ/gi71H3zw2+yoY+XSFn8GboOpsu2FBGIJsnCJT3nG82gG
IHWf0q14Mqhob5FXffQD8SLRpvsTWsgAW5zWSGfwp9DsFwzRtjrflP6Q+r4TPrus
hC1EC/9thhQQP2zZhBXJrQHhaK+h/Yy3AecNM7VPj9hwFx6w82h8PR3BI1chg3ht
PJuT7x+OBUZO43RSzIoHRQyrVBV/BJAXwpZbwyxQEeqQqHmvhKQJpiPpBAV7cNQ5
1FrHXLAglP0BwNhWlATDDlbSSjVa6HdtiCNYKijowESxuQWXsOqcjjSprNBvsNEI
z58Smx1uZL+3xYg0Rv9nev37yQUwx1Zfuf55lNDwQguRly/56nlRql8pL/FoVmC7
7RF1wh7ZYEDmkBx3GW1gekHKVdluyuTGVkty7Hu/abmgiXF9XZFViMKruVTb9zN7
sUIGubZJtN1UGuwcQOGfELOCEQ7tP2ojsDdeAlSF4xvMdWu34QWFHVAa/7H61XFK
mHw5BW4WTJsyJni28Dixyo60ve/khLg4huDvJZc6qmk+al5yfz5Gb62Ukksr0szu
KylC4kR8sdqNvBx/NSIxfEqwoHCBhCe0kWrBKqycdUlkM/7ckQYXHpeVhQY5zFPg
rg0XZ68OIhfhtTIusEPWQovnhoba4yEQ2ZQtA8eR1CQHaygQuZMc3xuPeuQfaLyM
8ABNIVtDSbTx+kfCQuHsIY+BB/QlUO0Z13ofYtlT77Rl2usVh+2BcwWL3WbyxAVG
FRJ9lk1bAIBX+WJeruiziID5UgU8tfHZaabUKy8cj9aJ/XXAbaQ3rMLP7TuLjR6c
KUEdqxkCk6QpH/EJhu7W8f8CEvAVXmRbyMh281mqe8lPL+IpmsbQs8OX+cKaAF4b
SjA0z3rLWT0q0Ro9VCny5Etgg+c57doMU+lHtVQwjjTk4vAQAVQXrFrBqPWzvJv3
EoCH/L7VnXaESVIG4D9esNAQ8PUEIcF3RbPbcpq9V77JF34s7ZjAWbYQdBMTfm+V
z5doarq8K58ALETIuerHIC2qZ4pwYsb0ZitqHTD8NYaAYxNc0cln+ziELx43hb6S
5CnesxKJcOhk/APIYyCbxfKTQxz6O3gt1Ic4Kga0rb4ZSQaAIDdh6UJMYalV1WV9
Kzz1Pos/F1QXQRqN8hhGkzQ/NCi17Y7pMK4DTHRAhhDop1J6r3uFZZsXgid2+ch8
y0Wy+9TESHFC6fShmp4kb+Emv1K845APlFKuMqW+nEltPCsLvPGQ3cOh9UAl8mFv
M5jmfdlzfDqR8TEtLHE03tpgNeUnJHrQfltR1oB821qcua0rbSuWNy3lG1otHWxn
dwFo7nYrGydE5vr8sdEgy9/lQNalTQR0fpmgK82N+mlrzxe+Rf4em32MNh2FS3La
Q9NQRKBawf/95eWb1tX4j0qfPR196eIOklpIW/CQn9I6OMzf3OAcVOCze0GDTQkh
q8SD0EZjpOEvJGSm16rcSr384jORbfL7gLcmpO+7pPL4C4joBmcM7dkVGjzuMpgW
mYDWCYaAgEp+iV0/w1SGSP7NsitBy2Gu8i0O8VC+UOIcornexhuWdKbIFpIT5fbE
Bb5NEZbcuI3xGLXN5b1KI5fbsMTiOzN9pqSDVLjeiwETkHuAYNWg2jjkVH+aI6jj
QVHbNquZrZ0S9qXJFfcClstu9WGmiWhex9jVxkMpuwK+OblzRishVwDqjS8viaAV
f6xYuaycLjkMXvrgz9WHQaMo0pMY9ESmrNFvfOgsy9gGWCwnC/b4mgGXEqt7+K7w
CqogSPjwQa39lwyuUiLA5MUTN2D591KoU8zQs72NIu2uUvDPGcN+nAizCm3MMGd0
UrV/J7hqaeToCQSF6N+k4fuB3Ax3Z5kDlLda4X2ZKjpffg8SzstrZrxLL37mqp2V
p9euMbCt4XrpAHzDizJTPDO8VtAWi4ayi4y+OWh1u6fdQtzYrruYUjHQLO2y001I
fsDY9PdbT5tB5C64p6UAdgxMZdLXsO2hZsQPum1NtiyLtsgzG9GUIBsiW7mlJ7y5
uqF9PGBW+9zoEbNy52ETshLq3/rZz+N6AYsKYjOkUCtAJpAYeJ8UCqVKmXYp8UKG
5HWm73vvEzJyH+FJ7B5CSnVPOAQjw62Dj3fTe2t++gKgDyycln9KLsYP/uQnCGBC
r9LKxF7VbWeX/bDkBo34S8k2kQzDo+1DKTBc5cgjW2hV+Dyjuh79v9epC5Ag8vEi
jpMVGG67D9SIX7TL3DTOkMx6I9ifgf9whDxJcMGB0lsdCp/ChOLTTua7RV0dgEgg
7UXM782ANW3iWHFmAL858sG+65K6+E0YmA6AE/z5foakJeVC0LG9hRHI6URruinz
wLRVl7n/z5gCaovQEQgp4COZ0jeD1syMOPSbW1XcwZDnuAug9j2WwTNx3N33zymu
9U99ojdxXyGskz1fEUg130EkocjghcRRTAiSiTQH2naaLo7+wrH70gJHMppwyyy0
IXUKbBv5iV+pakya1e6BKQxfOKXypcSsA4TBffShqKVpYZEXXwkjLqC+EDbQb2Su
sHwCtyFzXrlZkyh+1WSnApXtkPadk+pWivY+xxAitqXuzAVkzbY0sa2Y7Q7gk3aj
sa5lr4AOPutBsjmB0eu1ALSIE2+QJTHCzyVBRWWDm4GhiNxgWyQIOjEd55T8UOZY
+Z8jfivDch/Ki97QITVvRAyBB95EXKt/40ZCoz59lxCBuWrNZGE85HXwDVRexSKl
CqR5g/14Tf0urYLLAvrWoveeJQAZnH68kOULJ0ABL50NXJ3OUKNuc6Ep8uL4RRi6
q7UsrRhGFR3/xNtNJMHRmVS5opG3GrtmAewgoXQVQvNu1GYBv4Rf41B6nLaBaLDW
brec2qhT6lpYMy1ztjw96a1Oxd3x8omMZyHyZLa4yco5fHbpgeKNY0L+aYWnZM2I
ojtUbUSFdG6S98BA7aC7wwwadVUgy6bz/HNkXnI7hZVDGKmmdhcfg5xehAYLFQMx
ivDG7Oyc4GOhKpLogzjmyRFSIPWiOMDGCiB49zrDer99vZ5pmofnM4gyXj39ZIPK
0cbIpMkw8OmXikr58EM3qdt0CSNQruRuLgMA0SB1JzbXumkxhKF2qdbEhsHRVfRb
eKdMiVjvwOD3ge3jgKn5ftajNrW13P3tA6o5Zi2eKKKRkZ1OtCeThRGX+Uupk0Pa
Yswnf5YysuZG1npdsPoRxJqsWGDypPVxmFAExNavkUZI79QT/HzpAM4pcmHoX3aR
CzrNhRRnjbyPIM4NMVEXF+fTTw4D+zwoEDjoxexBUkGvbo2KRCZidKXvhMpOmyiv
nYlDFaegPCpYIL9AZVyXf7l84npHIztxh5i9nKKBZqfcb7y9gaXfMyUgUDZZ/XCw
cyWfeAKTKKTpo+4HzemRDezmr2YvIISq58RwZNp7CMQlB4TeOb3WYk0w3KuDub/k
hspBRVTYNUb+SOT43BjcyVNgjwE2jcdwFDHpxlH961Ujns3DV8OHOutpI0LVwevv
KAcraM0woH6XaqbI5QsqIB/7I896OP45M84PSXrMXqOULV2uBszvmX6xx7pnoWj1
R9kYSj9gz/f1UGsanazrUXd7fyNt0g/z4pVBrOcsGIQoI5arylhMmKTipjTqiWOt
sM/DhYEWYyhMy0wy0O6/HDoOOlsMKv0SOj5N1n0XBEh/Fz6yLoBXcz08NlaoXBE4
gEmXDI2ccmym1oTLC3ZbNw7M/wHNzh5z3pSB5OY1CM2fS7ShzsBGp8tnyJCMOjmH
5UV9bSkC51tx7SHqebFWbTxPddMz+j0UPK3nHbZ5cf3e/pLzZS1ADXsY733AbEG/
2tjbbRtTyqe564TH+/EzFjJFOs3U6aV9GyQvdEbneFOGngSzDutFDPHgEUiOmGJE
cOllA0DpSUnR7tmLsWogtOWAOAbsnfTjMv4eXFbaWSZq3Mn7tdTqkH0BbnHHwK1/
TE09VbptX/xTN8ig6tsejOf5ttY7J0kqY1E2Pu8ACMBi6rVedKjql9/a6LG+tWa1
aKN9h6Kw93oNSnzcX2RMkTaJs0wVU/P+w+II81z/6S1YI7YDft9i7UHriW0yRKm8
5JEdoYgfw3Xjq269+uisuUTLTMknpPu6zE0K6/4RLewqDqxc1ZPUxoZr8sJfTVoG
dAtdaaNI563DcW+GWXrlJh+eH2GfYkYCWln8mPm7Oob6KKFDr+eMy059G9WA95y/
LkRCfNqCZFhtJEb4aqiBizCeGKMXX0n+DgGWn8lSpjgezzIrZ/b+5564qWokLpjV
ffBTrXANleaY++3eveMPDhW+0trC7M9oawFPWT4iCClFN8sjQRj4tw7OWEgQAQLt
0ViDUUQFb7Ak5TMVAkngxeHS/HAeyoyt07cZAUexuhHIFd+DjkBVVq6zTxrtyGh6
QXPkIRo+Ui5o0APFlY0jCd/NT5K2IAkwZ+IGuUJey1bJg2VSrtidcOzOA105AGuc
jg9HfIR5WzCuJscX7ek/Qwtm5NPo7O2i8s/g6EfIz+6c0nwJV7ImFVuedtOGK7Qj
ifmCnn6Cr0NOo3UTmx77++/pEKMxIkLienk4EJO95ZuJ0bc5gUXLpBVCQQ4wgb6t
lG9+fYrkvexhwv27I3MjVm/u+WBhcsDM0pDSzHFTY93pGRHWW1N6giV1KECMs6Ov
DFApKd/GR6v5ybYMRr8KVnjxDj0364HUWUT5rwOiS6G94BCUYVAj6h6jZBk/MCvI
O3ZGfmpIbVQRCN5RIL9JACGXBH9vs71lU0G5FPMjP5l3OeP98fi5bFLt4jMMSA9Q
6zoZJSMBU3/AssdEKVdIwPVulYeteVfUuHTNdTzRPaZW/kOS6P7a6YwmvmVvyjhq
ViDhsiN+m2t9ObIyven57ANDEynTDrbxP5ADTZtiluANFXHLckBJOA4wHdNqM77d
FZCVYGvwmwgdy7ZSJtkfhNhvPAlL14ajzrH7/gMIVmAIkyZJoEFwEYyUv/kdZAAg
SLrxnMLEuoy8TRovOpPjG4XOA4mKHuSC0OUAWyvq0WrIG9WyRFdLKxx62Rbm1+VR
31R4TE3Tiq5pjaq1MfMm4Y8fe7ciAGcnNFgb98qnuGfrtMYdF80acVwU6SPIdWlK
rGInZMvldKC6UaCpFd55taQSnyZdahFeh3OAluQeSU8zMJ87g5GJCnPTqRRzKEcF
SWZkWCFhjy4+4+8Rt7goKZnG/6ZpsWGlfUhRd6wF73PNEpgkculL5gIxxzqXnvS3
lmMaLn889Gned4QU0HLXx4Os9IHbNJY19lnyAptZKF6tsTut6rkBC3itFC7T6kVU
8iDM+e/9TFbDLg+mraVDWgf9EZi68fySMUiCqbkf/YLw7yErlIRTCoVQY2VbEnkG
pk9/i4aspVFQoV+hpkAq+Qb8fb4HfVEVDWUq/p9d1U2fRPcMtzrXBztSyAwDUofU
5eJ2GmNmbjbp5kjrr6IqtZeCeY5/+Pd+dbuQYJBb/2Db+gXA399GfpLllZ/OEV3B
e7PiXrnMzLSQTquoJ5QnJwbCDe6Z85puf23m4gYkWDN65jxLvhM25R3q5s9gFHNq
DsfMyzZdLct8qe9CXVVzIktLKwzZH/M6/FGgWX5tmCxJftNYfLHNoc9gT6ly1H7q
DfVcB2XuBxnqJv41XAijtIXMfs/Dok88FojyvZ3Q9svWlJvVFl3JvEkX3hSlVS1P
Zr6S7cJmF96SyZ9BvqUYYwVDXab3DvqNasnKL8YhaVfrkrwS1VCY+PI8+KIuJwro
yx2Rrbk0IGmTr7zRreKNTMeklvGk1zxmrVzOTGkfCOq6GonBQVZmEiV4I5C8nrOh
S/D/4BjVWEHMCGVvDsN5Yi3WuWhHu5zo/lhy4PsN8BRgiIgkniCUZovqq+WJ+MxM
OBrM3YVEENw8vYypFzBY0THc7HEk0vvaMv0EEuLbrDuq93C7OdV6i13USO0JMujy
pGsjx0oHfFyRwnHm/e1+Pz2EzlCqx8KQPsmzx8PRk5z2WuKxNLjj+kCW6XzIoPeb
tFUBq1orJMdU+lb8Dx17zigE6RWmpYJkBen10wRaBkReCG5WSHTijvYOtwGU7dgO
nzav7QiNUA8ydbGj//qVD6AE03j6UFMoXX3W5MRaHZjTUA8Ay0YbONOFMbn0mGz9
3+4Gv5/CxII0edJF7t+6cjdbZAXyuvwQ7QeS2zm/+Nr+xm+5y0Dbdcl5V/ZYEg/v
zpCHYb0dB0JGxBEwEw9YBmDRiwAZJcgQeVHuaqQw73wHuBBAQFK2/s2LD73sTY0y
eAp8URu0LGB9TRe6+YzQvpZfwZ6+pU/pK/7m3a7E9c2ZetwSPuQOjk0x+YcNYZ3I
LyU2qp4FsoL5HfD9QTYQtQaFodeEzeQJMzUe2OpdYgkAqVucLSk6FQVgPbctsbUw
K8UOxG3bUS1LejfPl0ZNf0QcsL24g4Nhtbf/d+0iocC1zXnQun976vLqZGOqcodm
TSXvuuNrMQeOrCzlkOcwvLgYFeMjmY1tvAyDgW9ZIo6rRqHLeF7ytRy58lgmY1pz
U2POKTzACLP1Zib79j6GPPABGCEKi0DU7eZ+xd0ADmIuhq1hD4NOD4PrTycUddZt
A89ilRbrL5kRrdFyyAU/MzZw/FA+gxFKJCYksCyftp5LEXgfw4G2SqgFvTDPY5XG
d0Bb3hY817Bd5z6wzIxuhFAVIgpk/xsYiHbzCutzlZ/aaRoQaL47Y7dkZMe9NGRN
TQ0nDNAOBNmI0qDz2N7bE6YR4IExlyOE95N/iE/6VdQhhDFy7oAKETn4FYstaTrU
URUDyIb/EDdloVxR/5s5qBcXvFySB5rWLRz7vYRDz4ueIUZktl95b16KvKRchk2i
iwLooDJjO2y3kxtQdsZqxpasrsHaTsaIOijTyMXmXEj6N4nff7WciqgnbUx8jJQo
jNrzxYg8ZlOyBIeIn4U6WdQZb+xwXpB/QfqhRIyLysTT/wuM4ghCyt6UtLf1QuME
+HBXnXcISVqMZ2hiuytkl2PPYEIo5aFIE2VEknXhcU5QirxGbY57aJzcIYtBCjrV
3xs0xpbN+U7fo+qdzU5CdkpsVpoFVkbhjNZtFlKmuAsh8zqf3I7pVMzYLzqCsmHx
U6vhrdA5bIjgCCE+JZlzHw6QRB+wEI7N/Z90Ns7ao2ynlRvF59UX5c88TfpXLKjf
Zb5/xk19U7mrEVOJ6Af0y0BN4kbXpZ+KHcT5yxZQMHAkJ4sakfsuGeXfFAmGoVQx
CfZLIcfni9iGomLDisEKwWPYsDTtiaGk/ZjoVfxa1iQsgLltlQiuXisvqC144SL6
zMmj7QlRXSAFYLhuI0mDJVeo0oYCRMYqchQXsAOU+i1dA/o29R6BlzCS2bCjbwto
khhrdq6CpI1OeAx1aZKeLk2ywIn3ghqvY2IDMa6KFyl4KC1VXd3rtk1CKA0CWdjg
xGqfIKlRV3kdJUI88Vv2ZLldblsN5aIAmkXvMvzxEnIhuWOtyhAz+RE7oSMAYGCZ
EnXZgtQ3jgCXIGnKQM9k4KSZUMDdxVttbioajjpV/JFzTeEua+TahvWYKl4Ai1DF
7iGFq5qUJ1CMjVuYrkm8N0wOK/FcuvhdCpA7fbh4a8vz70sUJ2V4muEFk5p/WfwF
upzyEoMITCY/gSOuVI/olte/eGO2UlRRfxbBycbilCHa4WZn2OjJOSiEvcfrLPGS
hjtauir9NSQVI2rn7mIF1PRzOGtTQarhDWVbXm/hRVN8+nI7q4Wzi7lH+Mks/ISE
5LOtyqHyim/zVJwM6hjN13peEYjnpRF5rkIk0gL3WIFwn6pmagy/rMoi9vxuttog
ctyoSuk6UTQrS2KXtUEefQ+Zd4ow+aEx8RyzTiUfdZ3arP+HaSMJVGdI/Z2cGNcd
O0KUqClgVTd48QzVpzIk9pDpIQSYrdk82cAclO3mO/Ka7vuv2ISQLS2O02BXuyAI
SsUC5SJ7uHm3GqzwpKt+IGXLS4Nw/cVFD3bpLDTe9DCEdfY8x6uHN6Y4uHkHSrTk
u3J7MWNIdjlC32iIGlB7++ackNu+MVjO7AjzPCexndJn99/BuJSTAwII2da2WWYT
rJRAd/NlpIdCkER33iio6iFsqTlMF98ma9yDk8qH8Qycd8AmykfYPbxeF7CYmSMj
xbsCQKIDaiNvkGuRf14pB66rJUMmgjAWz42TcDhxGwd86Iu0eO+ZbvlvzpnN2qLn
oJDT8C96Zeoje5j387USKeVshohBllSymNMTBryv+a4yRTjmegl3WrFCuUo4Rjq3
bA7fMDB5S++tFe0hRBIvn3Q+9V6b9Ekrc/1gVsCyfEBSp4Rw/rgf56KKClR5Dv+/
EAKhRVR2cqo5YiyZ/iF6F9rj12zK+S71kwVz1QkXLhTKCNyH7GIbuqWncY+qj7i8
uno/S4xeq9j82XheLuKtoq7ZI69EgANJ2PDpEQIas2bPScYWqOltXNsF62NYv+IJ
keOO0WjQIXyeW9BiuwPAc9WRrUCRZkjTmcCs3RsICY+vR4kQIRfG36b0f/mO7QSU
Ks6QV0qI8iH8rbwUMxRsTCwwSRJ+Sbf33TqkZ9S1fVJd2mQR1n1fERk805b+Uf8W
IadY5QWSx0OX1SXiKN3NnlwV9cNa1TOy99MRqtq1tT+bU5N7S9DHFDj9JXMx6elT
DpYikb5TDg8StoIlzWsOyNUBNjadOcDvPP0xYXumyEuZMXI8cD9whvcJxg3QBMZ6
ItIShNCfNN1TZFr3McPzBEAMqBXgW5vH9XtPFSL5B8zzh57Dp3jC0KESoTYOWC6B
7Z7MJAnaEtAh0H1HjPtP8j38RKKlrtade4osb0mjDmntcYDwLqYryslKmdBuXZGa
qu5z8j7pZjqEoFCYr21zF/zon93aIo/qLwA79rEM2GqsOTiajcephtiLmWKUfhUb
E6T7wsswgh3uX2CChY6h7RBY96bN+N+OZm5RZsS5K+Ig+7filAUmI42uHNucbPji
c3GXXeSAMMhjZI8WZpAhQfmlvv0h/Qb+Ks8N++ybNqk7FVpqyqgqRc9bjbnQhXQS
19FANtgovqEgoA6NRVntQonOi7nlQ8RB8Bool4/LOt5BXf+t/9sXY3SIf5AwclyQ
brTrh9ABdUBPOSOyFEgr0T8BhHNCOVsx/K4AwZCpprhs7KPG6YVSeJSORHmFviAL
VG9+SxcOPUGjOo5G6Hy2RF8jsFgREWptzcEP+5iaJANqADn7b0ISBspAyQAL37Zf
KsJNoIEoe2cIiGTQAc/WFVyOIYU6vVTMa7ZfGfwrIhcwSs7R9xuGmRQu2LrpIuTG
AqbeG7Efwl2Mum6fC1vlAL367R2OWeh1nlFH3jIUl8Lkh7XVY5I/NVF+90pO5CUP
wh33tntQFYwGBP2LNhBRqJBRXuv35vrZZsD9xoml3xlkcu00YrPLuLEd50++tsrV
GsbFeQwudKU2EcUQ+xKxjjh/8vKKiIX3vpQyWzrtfd8BNYAfMwpNd65CqQ+a9MbM
3OOYPWW4BgZQsLjcARKbAE+cko0t3eXtGQOAv+mrpmF001No1V9iW+j1npWzjGTF
C+o2n+wPcepOXHnwTuQNN6DJzJP7ts42Jg4jxph1AS7t26PeZNboD+GPBd4CmrYR
/DeYqnjFUgXb6sksocSlqWZPxk2tYnvjW6t4dnGIJKzuW7k+JeLa5W2SN4jhAudT
ZTL5VtUz1P8JfIk6XPzldRHFy+q1V1mtFg0rp6P3u/OL6sD2Tr2sXkJUWxffumXC
/Gu81lEcj4lSRmS+6OvqNe6ERkq/yp9iqka1Ii+S0X7qpbc+roWD3Yuwp7SJ5XM4
NhWkRZlZ+36Wz/5TTPEATkOKvhhHEpK5EeRy+X8WY/OCEyQE0MyhG9OqcR7D0bd9
XuBn1822JNNFrN5GsOLUMWibpeRoceJ/eaxYV3e2u1E0TIcoxnNgVhAzSsQ9SEWu
bGZqd+gqUbGXkxiYhXDR6l4RQNguyTmCGqkujCaV7/uuXxRroPRrn7S7Psjxa6BR
9Lbchd2hOW5BXxgiDyvxif3VfAvPmY2XoqhrMR6fzBajkQp4VlOarcOV8nSoGhKW
9Tu+XR15SeZqulFcRIHEZCUkPkI05QVOdDmfW0TC1mkB0z2VmbAVdsDh6gOcPUH6
p6LLkd9pMGzdLl+E7/oM2oigo/3zajtLSTAmki4PHS1J4ngrIuPIVGcNneyLiHsj
LLdJkkTiQ8tbKMwRoUvlZKrsc3HMTOKG5MJOiY//c1SQRuh5GApGFlkEF91cGxEY
vbVAjSoMq1HbheIqJI7B7JqbaHzUhySYFRSD+O99dOtHNSVj2g3z+10ykmSKaZmf
HcEGQuTu/9+YHGjzHjxqCDKJlXiEcsT0G/yskkFcMrkrWSX+fpwtz1g5PDmKRCFy
Tk3y8QbTqaYIiF2THLef/iEjdbz97UMqiAorPayv+D18ZbfDYL/iokmSrQRDX8AZ
h4mISEZY9ZVLtqQNeo4GbT2oeU20JKeJrx/ruW4EOQPkDCYVTw8XGNpb93qjbFfb
xcyhWtsu0bTrAsl4PQWU4kSwD4iU6Y0W3ygbyaUScjmwR76uEgQ9NHrkGi7e7XbT
MyBk65fEnUTu7sf5vOi3YndoRY98NUZbtHHhyw/v/6+cV3weG5qndSf2G0+QESxc
BcVTQuB3r5XdktrApbng76pHrqnF/PxLMZ25GkNonJ1/rCq2OaUr3cjr2tjEK9aL
/zM7Kdh8oaHR0MK34MoM5/7IA6G9083NSuS5TfOkSr7VjrQemBof4v+psvINDrEe
wnXsFqf1OcxDTpYBWdBjHC8yF/82QDe5eXTz6EpJ7msLlNxjEl3doyeLvy4HjAG9
xuc1foAQCqPRgBVf+6+SB2kD34hOBFBQ9+YnGP+L04a7uE2OMBqNy7XmpViX34QW
IaXRjFSjUHiMKThe/vfDKj2xoazr0lj3inq83b2MVIxJXEusX/VyZSbt96OcVmp6
5RHAnRAsq7BpgjcFEJvMaUW6EuAd6ti7NbaezjNgQhpPbJwHEEuVY11QxcEPOBXI
GWsb/C76mrsKo3klXltTZ1TCSi2qBZ/7pKeY1wCJ+Bixtxy6X2LSqP35yx0mTGKz
a0BbolRqnzj5D+ggv0gk+jovRAe5PegivH9mBGqc/y+K59ziJcoEmW+BSaqxFdQN
PONYtrgGyjKXHtYWT9vt/37V97PUoGokZiHvkLEiiZpk+ckMwv7pEvPr8lgLklSm
l3ck9ZMyPg7dhSgthQMVDUkHuV999vHnDu3FmTAf7Sv4msxjcL7AJwJHpyxOf0VO
tux55tK1NEwj3aRubChY6pkbdAAfwSaXYUaVCiuKo47jAqrVOtFfItqp1/FgkADo
+T6qKMkTbTEtBhic5sudDktz+Dn78SyT5CY42rY0uXbxfU0tKhP7cCsTUhdaRh74
pTaHZ5vvS3zlQB+K123wnwj99utWBdglMsgNM2rFuWiXs+IF5WKtIOirWEsNp6y4
vSpfu/YEM6R7Z9DVEHQ5086MaVdCs6gLlCzYJC6vqS36iNYKoehPXBuNxvN8dUJe
Bjj/IQFai9Rpx6ZhUWJY5ng2U79HPHZab7e+xXcoOfBtEeiW0k8XNq6Vrbp8siB9
HY4cTMzy5+iVprnuUPkbDfow45kCFbf2UqzewHYku0eKuY9Zsu7OAk5eHMy0k9zr
S65TBIA3KAf8PrEdAL/18rvQ+hB9g5Kvm/nxsd4Sm+VyZexts+V3V+Gnan73kFHj
La6NmkR05BCn5GoNXNTqLj1zOSWTfwNadAOPSb/cd2iPcablQH4nuc8PvaMmuBq+
hdXSWfP3UHkn8L7vsMVnuDkXLZJ1tOEltOmKh9cA3TvGBrGMSv0woSizlWlf6K2K
EeJtAjRP45jabEY+I9VbDC5oakHRPCPGVRScZPoF3lvjrksYUWWLz/xe9q7ke0qr
vvDwMJ8T2bM71O3si4ud1PZuG8qyqk1PE7ppmjPr+lQS1nBUfOsz6I3WVhouzLcz
4XMZB/EdTMRQXsHW7Y01Yos4xqX+m/j9wPEy/opyy9v0ZPJ1eee/W3ISk6T4W0fv
s/VQKJBvgJbtt3SzUHWVvAng/7P+MnpDznjaxSi/0BU4yct/FEb27iuVAcjXS9b/
G4zg1AUO2gYFWeofu7MH1q9yxPqs0AiBRcCaevpca8TbaEwiXIofNooOLWPq/VIV
F4fOOIwh4lU3Pb/aQoofcNFnO2IT4jftnjJyo24MnYke6xyzfuVHHlmN35N/G9Nh
h0OKp3OgSInNT7zKafO732GM19Hxgwt1naM4wP/xadBalmWcjF1KKsndMRel7yu4
5iwHfRaNYPYcUjHF88p9rioKyDNBzvWVQgcuLOOWpy/JLao4fbiNif0KRaZY01io
evSOS4PqoqmuL7FszwCChr7Eb1mL8DJnMSvAPKjSqygQVOijRVm/fng7BjpHQNEF
9cGGrgDrciGZoUFEjSQHX1StSMiS+CmF52F7sTJBTVFCEtqW3htZEW91gWRGNMUU
pE/QOEmhFRm5Y7d2f7qYuwkPcbzq+obWvdQBXBeTLRPdthr5OPS3G6ggnBoGgGWs
KgPjloDDwNR+lqo0+ck30WIvS+9/1TRrhGbWdz7zb+2b4X/88WewhNtrTcRxM8P0
Y6LUZFy2djZ92VfXPbK7sBw21ptY8hm2x/+TPiqUMMcT+0a7VsF2gTGFgfyqHuoI
9IyfMIf+Lm9bQy9+uEHI8GnHZlRhV2yd89HwmAiyawxgVOlJd1qMAn2ivWy9lHhF
eR6+UlOHISIfyCcOkAqFFAw8lQLf/Xy/ocQ2Ma/P9sbLSLaffgtlLxkl/M1zgror
fmMHWqo5N2+x/nYS50cc0Mx7VPrvAgqIMTVvaRpwPqRmWZdVOnWFudcRmwl5CUrU
WZ7B2xubKu1ueJGCpSNl1FMU6PDKMNxB+J+LFGNu6hpkzSw8fUGQvzHPlq/GazFm
Iy6oscca1MRe9dkEe9t06khB4N5uA1u6RdtWg7L/cXsBSnq0WzZ5+ZYaxbwR2ztd
+qmLIPFa3kTHiuF966HaqJ02OlaKIpbRpZJ9ulMQ0972r/+bSxFlkW8H+tr/Shfu
wyXhka767mijzLxG+lyhOMrknEr4ZL0VWIPB3jgHRcyss0WfiGeoxJsHx7wd4tIY
wEFg2+CjwkcKMEtVplt2M6Tr0Dilw/NoDLXKVd+jqNd4l3bohhdDsAb2bqu4RVIj
00aTZVNj01ucCR90C2g8PnAM9oL+CCht6rBDZW3BS8S/E7fJ0+RhQe869dMs14fV
nU1oM7OYXzptgaLMJy1rkgmCurj9Reov7rEs1/Xoot11lAe8Kri1YT65fKCYNGs5
LeerHOluI6LwzDBbasTfGaLVHJ8mrOSOFBKS36Uu5FXJlyePOeKegxnXPY95K4Vn
kbg2qJ80HW8S3Vy/d9M8GvSFO8sFFDvn9grtOTGP7Qfa4hj37Ldy2aQEDuRoUPMx
iwNeapGx2NtJgzuaXJDm1RQlez2Omq1cUB5UbJaBH1KIvDWy08YMBPMtJyw1I3ul
5VB0Oj9CXerclProB46iardzOO10YTqgJuiu0QHhtJjlIEYbVJbWm3Kqz/8rITHB
djLDj6wfJ/fCZh/AXEdFhNY45SA3Z3mCOpAr17A5TPwqmG5O8plJYC+7VMGq5V+H
ySKQCAh2YwA0mmEVntYJP1jDvZRSPPlgSPGtwNXuFxn3FyhxU1Vw1oEz/5wURrE7
zkCIv9xw+z/HKeFMQllhKuiYEbk3GPTksU1RvR3b3QduF/rgqiwmIhQ5GWRCvOEo
Ks+sAvjRdlFdqHmblqU5aK4kQWiXMdj6iNGZND7raAz7wLv79JWXf1hPZ+Bd3POp
+hCMyzA/BRyRJB6sf7lR6sMtyHoutwQ+kTmxAVKiTCOJioSx7wwrzqmZczIwgru7
kK6982nXs4xh+NlaTcmbg+f5nhTClbq0HVR+FjQSOcpcOQRInthx8cnwEaxE7TrK
oyvNuvo7vtoaQA6GYIRZGIDOrY+yyUPqe4q+IP0Hkx+vQ8UXiXjPZZU7Q0Lx+F5R
YH54zKrsQh7TqwON5eIPQY3R1Vneize7qlUeyZC+D2t+6GkMYrf7mkCk6HYcDwVX
jdjKcFQuTC1SgGcCTVzeAvsQKUPg3AHgyw2aZ51sr7t7RA1V21iSlbFiGNflV4JM
p8/VEtRxMc78VcmVjKuiHOXGAuv1Y++D/9cMfqtP0ZcKiH6uB9QAU6wd29mojOM+
7o5Dgq8eYzqFIzmEXxZEAVc3GH5t5wxI8VM3OeYyYnEfK0G1ORY1y1Q7+XlNJkyc
eAxsNIbnnal6sdip1MGEwOCf/2YkDHUz+vxPwg6wBAVW0sxJXcmRacsOrDyyfX8Z
8oxYlmzs+U56L2E6Fr2jFBBj532agI4ctx3/JZoCO+kRyc5rM+4bXEdKDFR6odyu
XI5ooiTCt0yPOmjtC1hAgVRPb3/9/DDWBPQr64i3T43QZy2i+MRozqLlre9CfUIU
WmpgOk12FJnoqRKsGaAHP0ehXplOouncy2ZPwSlMowSk2IyFnMApXdU1O4+tRnnD
aLGm3OEIC8VuVs23ZJIoHaP2SsiS7Dm0+NqPlUW3xVuCJT80+kFpmlqQzUEfhNDY
3OIjyW2DQ89AnVNpT1Qpy2MdrRbzaVlCYweJcCnegOfZFOHfUDbRNNh41fJasPAd
y3MMTYhESeg558b8dT3ToJBhQgEOEv0cN3ykVZ5UPrD0FMCegmQMsHI2/rm6FQMa
TH5A9pu9ddWtOlr4YrtoAxSZRdXvs3tHV1L//ibL2hDo5KDRyOLSNnc781Xr66qM
aUfZ1N+Km1dshrzYKzuqJ6IrV8AZTS4BDXzW9BsvNb+APha0GGWPWKHG7GqNUc36
iRj/1D1cKKM6pTuOw/l3YyllzyrXqtRYRe2AJPFI9HO/K6UsDuZ15G6BprBON5HP
SYzZlqMCkGkfexSIzXouCAOYsRvlZP6Xsnoe3kC+w439fPDxDpWmsuI/yb/xe0Oa
BS7yrN8eoYwXjj+c8jqYxYEnb84L1T7X1ovgnL5QPXzZ1hsR+2fJ7QXeCwDv7nK6
aIjKmXaZGTQsEwdhaOq2Wl5/gjr1PD2HhxJyYj2WdQPNuvcOHgNXOr+OvRIyIj3M
EgN6FYwsKqxxiaGnG3YQrhR/VCnbTlLUu4yoMUfP++hdd3SSAnsVy8kRIAhYWWYm
Xe9q0w6NPsjCWJKafLi+nXOpH7CDDZf/FxDVwliY52YOeyZzwyDDTIccCjBXrfdk
kXhvhjLK84IHZ6Hxlf11+UKV1hzdg00iereG69wukW0NFySxUW9bTojopYk1sBE4
kn/TYYVbG+hFozDeZsVM93R6CXZwDAvuNN0mcQsw5cpfdO0cNfUHgH/1XxNZsw+G
+UebYV0YQpxWpF36R8Aaz5ba3XHsrhDw9gFx1GV1MZL0JdvGTemSWakKLsNPWH6z
aioORbg6p4+08//cai+elYrJMSVJR9T41Z0G2/JzPMcSsaWrqs0NoUNJWl6HADhe
iziJZk96VBg/r8mncSFk193cRRR8aXdVCf5+NdXtQVnIqjH8dviZQ8yFZyfXbyV5
UjHXhcGqIiljPd1IV2HPZU5FK78+O09V2RCE8td53/f8JbMiM8Nr3e+oIpFZA9g7
5ZdnwPnaM5v900JI6KQk64oMudK3rGtSMF8IZ+/WqfyXauVHRMTuh8Fv1z6saLJn
1LBPmOjdDzgsOdthDtF4FLp3bk2woQE+9LPeWjSvc3Ci4FWIVjKtXz9055I7ltJR
E3gA7qNAT7deYyVwrWKARC1T5Xc1p1c9xIgpuCOkpfKdJzzSBoHWASU5NayHGg36
FBcxMC9Fc9WHgsUTLngBbBXb+oJoVSt8V7an6ajxcpjkcfvdfR4QBaGd2arlzanO
3nXGLjyvsFb6dDE/IguATwi0UCpzoi/TFMELyfsLP9q/isG38CdZV1fpveylFgC8
YaMLtcGLH9sUgAhNs+KBAL+IPf4r3G3us4/ZQS3ZZEUYBTQ1tvmrdcdvWZWaYmSu
AYtgLvfPvathlv3/sqY8mdqWfqCQIKdlS8AbS+gwrWFbvcMDu8MzgNRKQvOlXemI
ZwHLFPUM77dzzAjyvZ613CqNSKgy90hAEScJOADGLifKXILVa0MaGnpslxaqSV9b
kxNuMOPJOt/vtX0wmvcN9aP5PFXKyxCRDQsNVgWIBedeDfVWPjPEQCAgAHadBKs6
99MGSGhOLeJgD64e50SeO3tuYg8opRvhkBQEdS3am10tTrg1lFL1JXzFCOPsAW+O
2D3Zv10VPIgjeXkeTkimDNo+Oj5mNWUDAyXNLVLxboEAOFhDLZTW/JpXDKBvIZ0M
5xU4BrLxpe5snMojBxEwqd6u8D7R4kuqvFVZDjyaYrRSuzRrCffzzzwIFLWRwKUy
iY2RATzyktRYz+oVQfAFLXbSVBejjiK7YRxL8Yesbl7IeDJUy2FPbEkNbT5mfTNY
RO3WcXzBWLTQ2L/RWSmPYNkKjaUPuK+jn/Nnz0De/SjA2/KR1ezFBhiCGZcHG4yX
qPVVd8TALBUIk9bgojHeRsBq014TyYMXnRYZ16H/I3vwfznLbO1HysHFdR29LrTf
aHVwiTESWnpGdHCtt7xOeu7YbbqDfyMAeJwshBCdJh1+i/5gytb5RO6bFkhcAHKC
pTwSU2dyne40e4atL3t8apRvT6BFohOW4VWXFZe1UT3/hNap8JVf2nFtnwvyunoY
8bh6RmHNvB4YTXlL56rYSlLg7CSp3DoJckOUTZ0xhLZjj2qR86EPyAF0ILkePFzd
sY2Xnx4NpmF8hg+k0xpk+f712ZIZ2WtpwdQpt43nBlvDs30Nx63xNFnEE3iOIZhJ
V2Oxhyk5cmYJwUAxY/xrn8x9jR1hRcuTUh2yc/HYVpDAvWoNBQR5sBRGy+qxqsGL
Cm7E8Z/mvy8ctyHBzB0UUVWw1ZbUrKPcBIh0ZJSDv0nXA87/OAOg2OlHQEzL4kAl
goEAzwpfvNq9/DfFPZ9DJVfXyzeici5e7ONTtBianBZ4f1q2nQF766gPLiPctHLN
TXxn3lAtNmTgGNC3j1FsaV3FTvCAq1f4PK+SJ/900f4iCGw3pueyaaTMqf/2BK7F
u8FJGcm4g0S0zUQ2qrKD0Vf8TV/0M00lOpmI60YeQaw1dgR08p6wKOBwM/5igoju
rTv4c2FKu9Ut5ROyW1kB9iE68BTxJXrdUcSEV7sjrUhfARQ0GpUkqyLTNbwy46bW
QmNN9u6z+4cQWXFUY+Qgo3iqx8lXOkh51hkAyT+2yxguFiutDh9r8c04ftQuWRU7
95vAAR7qyRBN9RR3wrjzzlj22deFcEBZN4vepQrkm57w4BGcmAgLs5dDslteoRXa
UM1uvLyI7l7KDoWqpHCtPy2PyYlDn8rohiHYCgKNt65oL7jh2Urc+4b0YjgqoVM5
5UGMstEWpuZS4V4i1ApSnoYEbytgkFWkV0zz5H8nHFkpGD5vQOQbWsuL5ZWomjnI
Uu8msGdJVokk/G6hBIWpkWTB22xCK4kuOxEIZYpYNPUCrrdYKwVtYw9GWYM1FR2R
Bq6bRO0D1IbH22pdta0gKEInkL3QZl2yPs+Qd+B2TdjzMVlVs1fudSEu1yyDZa+G
uITdAoZFC0X1VsLL/uQVQJ4LgSjjmt1cG7sytCSRbrFTM/l1BDAqB6Opsd1YarqM
6RRYdXo6KdZawT8mBjOSAqZxogJrHwdj+A8xY5mqV422yh7m/Jpd6hSjh0iDJ8Qj
jrB7rHyjmCccA4dsKCX3IajcSZqOKoHEDzP4zRiAITBGS8Sg67X9XSVVXEDw32ZB
DtX+vni/Th9J7W2UrOjRnHM14eBugGgMrjHhK3RDu+1KdtT1s9M15/60gLN4wJc9
tH8sysNg/38rFkWdAlih55rgxyeBJLMJCAb5cQV52Cq2E0c3OX72gILxIVsJK8tm
WH5uilHFyIBBldNZMjomE+GY95WaTu7toEQYkitm6kseXIRxfMVIkl1DGFGmTR8Z
ZYFujGOjQyxaWG6ieaG1XshAzvsdgnSFHc6bbwJk09BN6OEFTa9FZYfgFpifxbiG
AwXZHvGIqLL1CpVeA74CuDEq9f3g96pu9sGhAZY5Buunyb6Tvpf8u69H7YuOC+Hf
YbUz24Ue65VjXNRESPaG9bqbf1RYaqtNM1Rvb25iglD7gh3XlCJwOAwRhPgPaFRR
uCyODg5smkLV37rwryLa7ubQRLIqMq7uSwyDM4Xo/pNjzyIUWONgvFcyEXjrt2b3
lfCQSJ6Vj0yIsK8X/BF+JgU14jYJXVCKmgRWIidIzq6fusD8SWGCO5L4H5vPdt/i
vhrX7DUgOSPl7MgdcUn8N05EUFscy8HqhZ6ng1fMJaoTfZvDvJXzgRtyvvi3tPfx
nHXlgQ7UlxPlS6Ojx8nXqIVD9lGvj3sdq9X0IAki3dBX8aaUJzcrMp93sEpkeAok
oteYMWl+GZnqnocb4U5dXtq9F1wOQFibw0fvg4JKtF5mnXwlVP9n2K8+7x/23YwR
UAscMtSYxjLDOS52/971whQZKoztZeyBC4RTThbDoMX/YIQpUFauDdN8eVLA6hum
ZnL8N2/tNUBNYiDWzVXJ3Ee4whGKuii656OLV5b4FA2yS78In843Ctm8ENxsJQaS
mSqzpTKgDCUdAeW5KGT1cN5Ixqq01wUSZ+OdWIotyKV0q3Z8+wQwhH0RR9TH9cL6
a9T6CeUfUOVutqnjBUhQB9ustaCJUA+9Dag2BF14SHegYfxYESFMZff3lkOL20KM
6ynkYI8mc5/EZ9Z5xkI/6v3XgQmX3aoK7pQAlL6mk7yZPR9ZYqCNR500gSD5HYpO
xHccxzKLRV4wzCxoVHkaV34UP15NHUZtGYZ3dQP/FNMha13BJQ/ol1IoQgr7bhzc
8MtzPGH3f6JFT8wZ1tdCOkqX/5K9eLoLE6O9KbXUes0cH77IGXujYGsM/ExqOXAc
ArCvmoo4X7XuK+MK8w89YUmiZIrDct1apFSJSH3tyHWYsrCKwu4YAnAmCQ0VzZc7
JC1U4YsDF/XCuMrNEPCrDWL/gIAuwJxwsRuzRyFPIBGowjtu5D+7eBSh0KJjvmBT
Iq5wqNgqMaz21Gv0UvObxwd2uxffozLKQTXDb316w+X15j7H+yTJa6s94Ma9fO1c
xZL7xPIBQ68Wiz/ejnoaGRshf8JcsR4ofxRf+2XkX0hIRq9xrkLVADvPumrXvZBn
OU30IN3QYeGvL1GZqJbclRAX39EPmEuAaGS9hScxuDyDRL7ECnT5yowreUrimvC7
BhQfG1qnvxCrllBnMVBz1w+K+xMamhFoJZaEQFjuiGMK5eomrTreig5IiMZiQtg3
YiMjL6pvKQyZh8yWHiRH35lFdtFjkgnORo0iBOTgjbtu5O52HgDoaEJBkTG1Cfvv
QSO5tT2OeRUdF6SDZBJrDuuJfekHOzEotIxEG4WihQkhhkWkX9slGBKEdistgelz
znzudHhR4Qt+/y+5QDxD1WC/BljUl9Xu8YLUfOkohunbjJBF6/nPG3/F+yRFr8Kh
8bfGbVfYaZTji/Xu+DiqYJ9EdThMA98CpdZgzjN0vmiciHQgTf29yOoAYyHyUOWZ
e7YuVqsbmQe7SHRuBDRW7ImSn6HS1H002uaWs8dEHQ/kf1Hla96qp/mTzEsgTLgV
2mqRHVMKnqACmZK4L3TsGqmoxjruSEJ6RdXEm+jSQtco2DngdhAOKKUzeJpmx2AO
+VRDglmAA6EHuZVd10EG8FDHO/vIhs+bRlK4jr4BkGd6Kb0+BWS+KIphTu8nHgP2
/iTNauSbl7S7qpe/43dAO5VGtHt5S36nWcgRWFVlczRbu/sWA27Ox+16ayr2w+S9
TINY8hsNemBcmWZZiTJQdjwMJbhjUqFllHWf6cSI6Yk0+FqT/+ZqEAoXFl8+d8vy
c9NHYcp5tcyJfwM+SwB6noJzyjXZtXyA0PouiwoxDAw95yg0vdEMRkuK2taGNYT7
fIZYwx/BNSDvymZjkgdX8/o1ikjaF1s1Ig22dlrKwaYyo+Taufpf4nUtjlb5E4sz
TgFnKHfFvNCv3xqGgbatYPIRxLKdNQGyJ0tLbvM0s9iFc7fRV3XM09zvunh4Hdpv
nd04csIk/89VjJVMj82bYivw58M3NOy3g8lp0cYPBKZzDhzaoYyMQ4LoXSCLwOjn
NC8kwAOGkSS2MW3w/1FJxQaH48WPjfHGvVVL9hvIom6yESG2nAT8bEpr/ipBKAd9
/Eyhr0RWU5+80CwmzyeA13b2mzdiDmic+qbPZixY4ZCpIiB2wOQzEY5j52lYzN5Y
3owx6/SF7LGaTK2vmuVyaiHAfuV5PaRVpvE1fmnWZCxVh792mXm6SPa65oTV2v06
fdW+UAD2F0x5q84AiX9nMArsni/iWlAOrbQPcvwB/nNH1setEEuUo5T2a+2TXdzx
cgTNuCg2GzXo200+re6eKNUNATur4CQXavPCJW1wDPYnuLs+h8haQRgU07LZ2Weg
Fo5D6tcGqeeeQTu36SyhAzCwwHj7iQ0gxSFeJNYWKMIyZInQdEOsrHrMsAGX0rnI
zwrVM1U4i2QcKgNUEUa7pOsUarSHA3VsE81WmJKNvjYFzRWPlrwzq+IbdG5XFK1F
VMT6LFZpA99M0y66IKWAIm8SccgUBVXkFq6vFjivy2Sg7ytNXS31F5qeFt+N6Jv7
UM4zNTef9TDNP0l/tVC4WjWe3npAAdcfEx3mGez5MXQ0MRlfqZ4HVIDXCQwlr5Dw
nT+xvx18h6EjkXnXOVx2hvN71hZyWhnVupEyLgVo/7UXeARjzBuml0KelKEc64XE
8GdffrDcencZct0Ag0oJB9NMzC5Gyzk0ZNWiIvgOSKBe4XT3tE9F2UIad+8b/SqE
897mfBFZAF8JkhXlLUBzJed/a+IGuLITAC66KuL3qmuZrr+GhN3hkRPmhvuk17of
jZHwxawnV8yg0KIuwT3zk26Mb0uELM7lfLED4K4OBDxlIL8v7b3AXddGg2hTQedi
ebb77W2lNOpZxuqigNZNstcyox2Y+7D/5yco5Cgu6giUb5PDSmCCq9pTkrp3iWKB
0IYj5dgONvdbm65o2ZEHBE/JFDneD6n4PiLGIkJN+UIdW/JGmsatLduICWazHie5
h3W6Dnuq4KXtTVK7u3Z94PVkdFt/zXZcf/cHqERNC00KhpD3CeZAKkhwZYsfRJq+
zdz2JHCyAf7hXvLYFfPKgdu7x2WnFT6j14M95NOnsWcpn5y18K/RIV9FoxvJMGDy
cl+4BZKcAmWbHlcFj8LYdmMx+CT8nxFMKHYd4lOae5Sh7eRWrP1OyhVDE06hw6QT
t6mJlY/i82W1kSoSugGNl+4xZ/kWOjTrmNFDzVe5IephY5mGc6mpizw1gc/JLDOk
YCb7VamC/5PI5kToSX6Z7ETzGnuvAMUfcWwTFmxHBvsiNwSxpF8rnzdUVzOk4i/L
Agj1lBNVQpEcoLGoZfpXLfW43R0n2TbANBNCCcZcV5sge/LM60xOzAAmA2MFZ+IT
rMs0BluG+v2DALwGZvZ0uCGXVUfvH5ez64BV68SnZlmrc2wzduHTum4LpHwvIq1E
gnHJaUGFj0ID7fzO0/yG9/rQvmBGG0lx0+DUpNQbUJYXCg//apWg4E/mwt4e8z7I
Svra37nZ7lWwRoHvz0I3YxHLN8cYhNKZ7dtmGp3LWGFGgVsT9kiFh7bNqjvHX8rU
nI5VfqY3QYb1z0lyJC2rmATw4KwOrTOJiHjEB9cqfxqMq6AeVpv7dFky/p+Nt65v
wYQ5Zm7UPDAgPKje7c3Jm4JSGiSDjXq7hV0kpZKmsf9nFkXEusBVqKyIfKr2CQj3
AnwA1/seJnnBpmeg3jQL4emWncCNyWN0Jz4AsTe9CSrkDyMVDeGtQlzPc/Aa1NGq
I3l7b0osVDioTd+L0lK6rOFaCLBH3xjiBa0tI6bQzgtxyqKDUfLlH5lVCInYM5Pp
AhUM3ZAfyeGjugKsH6ICffEEMbomeJXQxFmAZ2Nq6bKr2PJiqyRvKyk3hjM62Clr
WWcBNknX9IBZKqj539bZibhSXV9N/DTrW+OanvkMLsX3PA5Oho2j4Y7UftMPkeT+
4WA1/y4u+KJLwv9ANcS1HR+9qhHgKwHxslHYcBPAQLclLn+hy2et2ZyM04zffXgg
iugXZnl2JZOi/LG15pbz973p2Yy5P3BLPdd6vZtPGSmvHPSPrMekB+R4MJT53om8
aR5ALMuyzhFzvrMtxmzIVfaYaAz2DqWwkKdU/SOnNaMaXoxpEI0ujkQIafeAYNT3
rthvCybrF2niiNiyzeO+6NttM8IGIVZ08kgWnvUHg20dVcLdYDxu8czup1DgSRQ9
7VTgicsHe73gvNpeK5IZVnTw259tZFwj6a6KBhCJJrSOtPSImVm9kDjqa7Xum/QX
8aJO31fvXGt+amunpHikY7UALAJHymuZ2UweJb98nMjdu1j2oKLnNGIGleA2jM7X
p/lQrmkJ8DdTZaRI85zqKYrkahSt5AyCxUOi6LX9eQiJ2Mk1JMBKtZXp707f2e9f
EAknfY7pofAd5LZieleA8XMV/ODxiyEi9DiropCbm62wa3T+7OMJBYK/24BoUz8Y
rWN1zHnsVgA2CAQ2KtpDi0lBU8QQLmE5xWH/4+QA6NWGvw6ZM6X1NcEXOF3XG1kU
HkNi2Rancxow3NVEU/5X7KBZbf+X8+tJv47uuQEkoTuphOCAUkP+R2F/PkbCHkq6
Now0GwiN6s75coFbJxyFd/YntgqKt0/rmiAqKwpiPay+IyzocDS9esiGE+lA7t6E
W8NSQuqQjiJ+d1HhxADr6Va3JS8oB8wwWJa+Y0Ahi8iLaZiNSZlFvreLRm2AkKOj
t07P9+AItgaPFoHFEy4vyehnNVCgoPwXA40b3aEUZHkbSCavel9lwsDSXsvMBKcC
pXOnNEB1tYGZh7RiDKRBJBidlse0RzcBuyXG+3lrLWlDwtuwHtozRUy4cQZDZYgY
cd8Vik0lEUyWIIzaMEMw8iqPUuzTey23Y1wjZgg339esVv7BlDQuFJ7Xl1Nd+fBm
tLtngAyn0jiAyduZYCOOTXvdcQHPakxTAvBUoaZ7OZuHQMqrxi8sM2V1lGrjksEy
X/ccadZaEL+4MsVlb+zNfEQAHFltFuMzkw6DYqbqPg+OVRovILUwSur+LOExyP4a
LXgvm6S16WBVkK4nyM8ZoZe7clrjlG+bmpq+Pa20jEA6REW0VUzAfrnwplOEqmvW
21TygQec2SoSEq8eqzlX9Kx83fgvZNOwK7Zxud/aswlTz1+aEa0KYfz81ujwPbVu
FuMf8LMKuUcL5YudT6B/I3GmTG3kj+esAeJ5bYAMNZ4OwdDZgO1tEmE790/sNy4Y
Fj5JCuFmelfiPREc6v8ES0DZtPh2Tn25vUDli1ic/Sxgv9QNNvsYizMbz8M1M6UM
A7Bxl7CAqcXkY+atoP2GuwicADlrCrm83oScxS+WdPFBC4n++7O63BXrv6RkEAY5
5wU5AfO9J1RrVYbkXRQEZX8BydDfq3dbuUZa+mpLvERKB/cZl6OD8x9Lz2IsXEmx
orxpDE8kRQ/niYr9w6GirBW8hfjgrKuQDmp56+hcrEnBYm/dbSag7NHACkBES13b
c8KdB+C2Uf7eclS6T0wdRdLt/BNVlPLI1kg8Iqnl1wgGCnk3ksMBxTkXX59uAWWu
PoEgQJW76ZWtdRUZnOcNnnNEnGLwPgtcnKZcuI520z/rt4XJCsdlfd5X3QMS8GTs
IWWNR5+NW8XMSVlf2ipeNa1bQl7FH4pnJdhxVlZZ5oGy45x4/gVfh1tgb9ETSWxa
WyKgROZML3gfBGW2qDkJsH8a49H7MpoZhrV6aG3UUIiXaQcyOaslZfjdllc+9nmZ
UR4MCPC/crqCnfcgAYD5WDQsDhGPvzx8dI4trKlkfAMVAqKcRvLaSqc+gEGi/iRU
LkKJbD+PpQ6VbUnEaoxKon/ki7Hlosw3HdIrZXIfLhn3OhgGGBMf2Tz2UxPwSfLY
zKT9POxdGxSP42fjiW/RikkdQbjPE10SbXPoVrZvVSHq4GykybIqepZl+A9sUHIb
W87TppQoLMt5kPZaQA9iP87VjzbZOVSdL6OlML7z8dPXgW2E3ZesFhMGVhVuNdaY
SAjtN7bYwqL3onOmN1Hz2ABuTTWc/3LuxLtksbk5AXRFK0MjVUMSm0Wso3Y75LvF
+svuyqdtfLnxqjITu6q/oMV+qzi826Qo7UjtxOYui+0zBnhCs/VM3YhzN4NeOfCg
1xdEjrhNIsDiPfyaWMpjfv1l5deKNrnJLBw3mbFesP7A3ifyr5GrhnxoPxF6vho+
TrrQv3Y3pKc5WuqzM3el2IGGcFG46ri2qifZA3CLIAPydCNMnaHqpfR/x2V4kwVs
qO+uMNY5XXTIxvQK7Lbd5aLauZBvl2/JN43qJ7rBibwdZ36n0OVjhvc7Zr0qTJJo
nQgZEuGfE6AIdFtYsyHUa3fDuMUK2ZCNStCCFhNVE4W5v7ilmV8G8htjlk5KIHoR
eRn2yWQV5ZwagZZ97OfVqavvoabEcWvy4P7dOz+eMAPlJBo8gVjNlO/RDprrvhOJ
iCfn9zmDn00756hEPd8eC4J3SsIMBnm5wqDyZ0ySJ56/9QPd/h/X3pB+njjkbctg
f/QpObF9g7qgPBsJVlrWPtO1XHNUTil/495wMsuh7N+xuArYegASimhWuTIymOuL
0QAPKV5RjP7KZKNRcyJELDue/JWVDavwZDXpQKPx56Owakns9saTU/XPJpQCDMMp
TBzbUjYk+M+55JvCqf32D+sD685CLvJ55GEgd3cn5SRU2/Odnj0K7y1rjFIJv+6G
jymaJZhteXj2pD7tu60qp9YcuPLdLmSbL0g0BueEo6dbTM5vrITm77D152W0FqHE
CN3VD01kvwmV66oXZVeBcH/fXiNn4AuYh5i3LMJwEwKmHF+K1imhBcR8OkWFZB4I
wDvZqhlvXSDCb6w8CfiVIuJLzwt0fqCFBwd4/Cl1EwseDJ/3oVsIjfArfaz9rU7T
GGf80CydW8UmM10I5u9teybwOxr3/fSOb9m0aSHzUE3DkURiKYlG/AaxUVIKCO1W
GSt9nWg+8CBpg1MUeY2t6przTlkzPiZirCAY1rfv53hoxZ12S71k4qYeUyAZKdvd
QdgRYElKBUEUXJJS1gjFhEKXkJcshZXJ0Xjo75Rzfd38p21GHCP8QyhPzIqjAKoR
PLViS2B5tP6WBjW+LqBKCFvf//lCtHsQ+gfZI3IfkU6jDSYAm0TaCK8ErFA0zyye
pdA3bsILfjGQWYiYui25pddbmm81U4ScNQQft13UGwKC+LgXiY/qw1pFjYEkz5jJ
MTKfuEjcyKqQxsiHjgshwErOpbbyN4TsNkNW933FSmOxgXWq0iYI0xzLbycaGTwR
BiMO8nMAvcW6FgnQKIp6rnynybT7+JkVzoe19UPQcpw0UAq+xe5MgGCJj+2+hjWa
A2O9hxwGlKwApvXFySypOy9t+O33xyoeNQHk5T4Vkzx6MViLjKilBfB3y2/R2Zcd
Gwgctbsi8IE5STT1xvvjcNatmjdCQ2o+bIme7G6wCuxqAbIYMNg0iqaHl4uP/HuH
nRKFGrLtCvMB4xkoEWSZ+3s/CJpyBnSkxQwHvPnXvyo3/uPAOP74hTq+tESIUaio
dyoVLZu7+nFj9KISWIJi6IAFED5GODPGmQoh8HQLTNTsjK+b/da3ikpynKcMPiqZ
vCv/Sw6FytPiy9EqcexTlPWcYBZNsg3Xoe2idc6iBUGN5uRw5Kk8oqoTHQo2iq9p
s0zRj4o2LJeF1EViF/XpyT7iKvoL8NoNYf8hW7CvhBMQA7w7uwp0Amr3VqMRD/Fw
3VhavbnzhCsztMW52v11u5+o0tbgf11nwaDL9UhReqKI1rDqjkDEjG/ujG7UPDlr
opgGqO/z5btIBG+0IeVXMBlvTrNMroPTvf5lHhmMDVvU+TfP3ijrPmnPLOIGvkl2
DFfdkgv/Axe2JZJLrZHAGVUl8soO0tNvxlH+RKqK5eipDR9hzYUt3tCZEOPp6NXu
h2+nI5ClWcjJKs0YErKgjFbX8uwWJtRuXMvOSAy7UtwgELxKKuOKrXMTBbgyzB1Y
8EBqqsQ81ycVfutaNElK+gch0FZ24K2OIPv8GCbqLHNG+J6u4T28QtGDhQt2YZi8
BSBQ8zrUBvEesC8PygdMXfbryCA58KvAGAnzWV6BPhjpN0oom+8R12vPcLkr0mxB
yKHAbUSm/tgkEe46k0FmEoyl7fY2W158jyiD63zNNFQRKFO8spFGauiNMW7ePfKZ
Z6YLxjY9sSkNckd4PQMjBSLVk3JCKaMIWMO7wOcdhJKngXV0mA5kzfeigG4LAyeq
Nt+5oLrbD7K0x1oLoJXBUQ6TBJikjnRKjBdrMuZNqNY7yCYKH0SnHQj5rUBNU3ZW
guJMkKAClWN4qnZLlrt1fPkcqzWnODtyFZ9si5YQKSiyS52m1b1dAMlCsIsb7R2C
hl1WGPJ572BVWRADcNlM9nKIDW+zibVERjGFcs83ljvRUvcuMAEE7KShvKymgm+V
tDN5ExVolaNVs8U6OpGuFMr15Y1+3qHICSgg23gHUGo/CtgjToGW/X8RbXvNL9Al
TkuTH5RUYKlhSenUKBhrr/GmzPdfvZ12J004fJX7HyUyZDllK8DiAqZPhH3Wbl92
ZEsc/Y5XUOgxDvp2YgPxXScrDutRM7tLPNdwhptQNgDhXcOmRUQqziqfX/GAW4lP
NQtBUkiTTN7S6H5gr8Lw9zAvj/tZcOTzoDLQzlvFBN6FvOmgAaomXNFlGIhGho6o
DhdBkyDrmw42x1ad7DpyH3r7jdaSCCxum0MpshuZabntfPpnHBQL9oovVAW5ZGh/
8MqAQGrxV3iSqd6UB0r5DK3urcgCt8hIdZV5zAYf1lsjlEouU1QzMJTRDfXEq29S
mQiJ4coiQiHFAufQ1TPtRFvAOOtMaVA5+If8yIGcsMKZJBOTiP+JxaVSaamtPuRs
e2WBiVdq750VfVHXO5B0olBtb/TTM8wmtlzln29zDHQlrRG08pRSyi4X63el3Ezw
FHcMDMYAM//BCrUU8rOcJZqaCpGeVFny9BjSERXD07bpRRIA9Hkgt1dXEm2Gr/P/
gFpc7Y6vkdtS2Hf9A0gKDR9Y8UQ9H5orZ/Yw/X5h3ruqKisMqgpZwPzt2x9Onkkw
5A9kUg6ndHjfB+zlNnVfc9bk3odDhRl6rSWpMMuWas2bTvq0BFH/U2dMN495Z/fC
srvOi2yqQu/HPJZ83adi59RBNG9R58SINpz/hxxL+D9g2FMBmdCGsb9063dtHFzD
XVGzJIZPC607egJtAtGNvb4j50jcgLEdB3goNPuUygwYnp1XwfzZkPVoycBvRV30
1o92uEX0MS2Zo3XHC3tTm8kuD5taUOCyKjVCPdWxGtl+D8tdfA7FH7ZJ/ahxMpDN
RudPnvk7kTxHWGP9nOsC9ldH99uehqcr4oW/1qu++fs0MejZgqtgJUM+rV2TvTr3
nj5WE3HZCmq8p9frFKJf6ZZPNh0CMGdncdmBpzx39sujxUz6uJD/wHoGcw0XVV+L
B5kstb+KC9Na2rl0v+HhCV0ItE1Nq0vg3hRFe9N1wTb3wAHrZFsMZuXfd1UU/kod
eoQQzzis1w3z4hrr9FuWWgoE5/ZIzzLjkf3c7jrFVZnXXN5bJTX97444J8iEitBb
KAL+vQLIdgXW30+b5GOtJnL8m7KykJHaPrODVpmbMkPDE6R3FRxuSmqhV3g6RB1m
ID4e0JRIRKIvZqu0x27OK0bys1E3U1avqsCGuaJTk+XUo6210JmCwtRd/Wj1bd9c
v7/d8LAz3Vhbxaw4is7hgACxhzGi/IX4cq113B9vDHcGjR83ChRkj/D9iX9ydHV6
snSG0d/sCmQPpIsXI1UDpdAkyEMEd/2Rne0yyPB2XwQiO+xK+GFO7S/TWCbYIjdF
WAipQpu76ksb5QuO/7fFOQiBmPxA/Ons5plMnmhYEPfnuYDfaBw60AdVefGa4gvA
c5r2lQ57C6SZ4E9M+WmuB1SPQDJNkOh4WFOrZ/0kUnvEAclegvqFrq7GpMqQWB2T
r5MUyzo898x04opoggZnRjUNfz2Gigy8DsHv3gsCqYMeB/obXLr0KIe5pwl2ENW4
QtSWjLXacN6zR61m7MpWxirM9a/XbrRLq/ced9lsAMb6UwBiC/4NdFFKOIHlbVln
gpamN3lxaBt6kPwbfdqvkaRa+3rk1IrBZcs8+XuXyAtfXt2CEOUADHOsfP6YvkOr
IB0SJnDF8CbnedUEj/JIVsB3cZdUjsFGhrgbrjA6KYGKcV2qPkndh5heIWWOzg5C
tlbUZjFLyr92JcXj2wXWgFWZ0QTLbeNw5LQLt75SlIxUhBc/mMtw9ziWwN5GPEuM
v+IUI2pHN21TCPSG961DZyYAgd568MM6kIWASSHHlQsQ6VAW8PjJJjJELnEQ9WAf
/utG2MPQMS8A+ov7XTCTo7emLqMJ3w3KTou3GOn0KYhmPQ2OdBpSCgCSMd2+0EOf
F6mfE1XmW8hW2oJl0VxiS6XPHtCXdryXrikc/8ZSKRp5ptdLiRcP5f2KEEEO+CS8
DpHQtpAmqZ5SV36n/m7ielKY48YvzJBMRhq81KGLlvXIMtdl0lBNeAzo3P+zfUAs
`protect end_protected