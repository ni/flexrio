`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9056 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
DcaI24013a1ntsbbicG8fzxP/AelpFJgvCejxNWqHJdC7fsYESvx/K7Llpx4eaWA
X13QGIJ+HbosXQjadlRV+6so6KilJA2JKdXSyP6zzSvoRbgUxOhP/vvGZDwFhfRf
iHt0KtckNppk/L6du/3i4JdJoDCacH80ZQRivcH8EY1ODjd5Se+kf4pHuzZ9tZQo
jOkLfQZ0O4w92NhjDcBAzftvMro92+xFNszFX3xjTF8Z9Mvtfx+US9LEGt+FznCO
hZgy2OD2WNA1RmVsPdlg3jsffFgLTbN22K++U6Ovx7uC+liHj2nLGj/cbw9o5XwL
ofuuyM0WYzoBejOu50pFli307Pe+vJhNfIF1p6FJEcMfJilPLEKE3M0VJMEMLRK9
WFv9KFzO+M3HgW8xnmVTN2e6pcOCQAC0GQcSg6DkRHKUokbFiodBHT2d9ks8WoK3
Xrj/JT9UEQ6+c5ha3+HUQLdJKScI56HoLYUWKSDlb3TaWuffooSWLjDdsCkg/JbM
O9RbXdousYpUHEAGtbIECHl6mGSRWi+HsICWFnZMx4EAsw909CE1sR3mry3BjmHX
COgD94CEKxYHieHmQ1lrp4wFQv1BcfJbARs0gQqcQn67FAlLYpE0FJMavS7C+HH1
USTL7MV0bXzDWuxlFEC4zqztdfcmeNXGg9Qd8rhqFVIpDuLKDT9KgbLMzfB1ZwmG
jagqU/hY05dEFvKHtZK8/2HO3Vw+zoKrfjsA1rcnIzzVh9lHNNJHounCzSSlC1IY
N1QMeY87UVVdJwidkgIbSd4jS55NaREyurFe41zq8LE4qoCZmwFJAiPxBXv+jTXc
sq0F59clS9HTtqRVgVlNzQiqnKBnnxweAZhm+rJL05gU1R7Ytj4sfjQhRyWtOs6R
rZRbSmcYgLZqsL49Hwj/gtchBeZgfoQSrafaxqLMubc3ZWyEVY2FAgbcg9YWO41u
y4KXp+Cn2RfYn92hgSQp4VewOembf2BX79AARqI00MCwVT0CmIeBahoCg8KRJRKb
KJxv+D3/IxMEa0yPUHd9PzsiGUWquPd2vysZDkFnyjK0BiYJl1FzQo/cu1e/Q0EV
9wQTHiqgv6i/3hvQyfHB0zV7HFV4YF23JfKArDJr0rgxYI5XwJpD5TRfc7x2Ay7W
orHJlhhGmB9eF8ZvfPSPm829xptr+HST9u1ezIab/IX/Q5CfZ41crBrM3BwVVeT7
OlmTgez5dXPwgffbm7LPZdANB0qPH2PPFcCkriyPlXJ5oPQ/c7CeFxUS+0fHLFFJ
lDz7MEKWweZseA55wS4S9OcUti5973OmIRzHSHYCzhmIQzujCiUxkGOZc4L3Iv0V
g227yUKPMdv1FKlJIHW/B4PrBVjiaztAdLuONKxOk1lieVa3xTCUIr4cfXKjBiye
pcrlCDgMVeTpIvk9jAAeSyyC7rHdgsRn0RybrNuseT0zpXeQMvF9jvq2ioi2JpcG
9iUwFdAg8QxpHLbfz77AriQYqHjwmkCH2RXJ+0oeK+HmgEvj5dw9Z8XgebbSNFWH
7itHxlbEGvHA08IJiEWg7sCA+8hVX6qOGssrHjJ2xJTu2nYpu/j8YzjS1ZMdTsYW
bGASwVcPQbjU54/bwg+J0oBxw2VE/luBHSPxkefNA4Hzth1ahC3xaY3Ku3+Nk21m
dDJKc3NyV6no4fdEib05PKJA5m7BvuDNctTKn1z4owmIG5sYHBXereSc9WEpBhtG
LQA63jkwbEHVTXjKb13zkdIvt4JfNJARtXfIH0fLPKhavoH9WyOX09+JFrekgMay
bIkYtLDlBkpzoNv4hSyRToQIc4/bpaM94fYNik5slrVhm45KWdExQb9T1m0GaKac
KMwam2az+eOSvQBnGmv+9/igAx2byemmGoO5pj9M7okcpXT9U9Ois7j+PgimuyJK
H4v4N1XwomM2TkLghm73m0bsq4JHZ0igfj41N5kX2lOpOmnH0GVIpfeHWnz9gCaP
vKO3oYAv+Zh9yw55gwFxN5+Sm5IJNrCcScNJFaf5H+A/zgo5014ftWp7lPXJN3ax
CS2AP6mNxNJpwtt9x6Dmh1Uu0pLiTVkvludZTnW90NfpUE5VWO2ErsKFwoXsX+WD
xemecJtmQAwsRcDzzh2Tv2MqnXpF+PuvfxemDhZfwuO8jz3U64TKfP2atXtWN1h7
hYtrdYsCh2Xix/M7uSrgKcBhDsz3owt7ctkLKsqg+iJfJsh0Qy4cdNQve2ftfa8o
zFBk8p2gI5FNMGaOL3IFHIYphsO4Wo5WJZkDfsLfI8umo+zNozjTpeKj5tfZYsXd
43harC+3h7mNkscd/3TEIeIyc+IlxVss30Rx+GHBDwpyUyVnpbGsfTayI7je3JjV
WuUPFZL8oiMQoR9tEyUBVtZxFD0N4f5EMXyvfYKXBzSXtwt3yu2+HEPYluuqP+xQ
AqrNvMYXQ6USrzJQSkGtKo/ONLj3175iyw311uHEu6NkWAoBXAf/gP0DrReEy33n
yQS6mAiw3FRcJAQ+ZRopF4FWx33pjw6tJB2P1HQ6tgn+g9UbHcnXtddzqRnGzXx+
LPCcsQGoFCGR6uXIY5CsWHoV7BWd+x2kqJrEhBQ/cdO9K0QOCw2lh6vKXT4z07eh
J75bCmK04gNrxNH3i8t+w7Y6v5Z8xAZNuqDuZPtgaf9MvACr2j7vFJaGyztazMBu
8TLKCbGYMkeqdeQGqggU2/lIOc1EWvMAoyesHRr7OVuoHfW79g9xTiC/KK5NlWO5
P2PsS3JRloRbvDfgAUcMxObfUqjEWEpSkWjVshxKtie5Zi8xu+ROg6Uu3ZUyLSUP
mZEK5V2zDVVGI4476rHx2MaRrftK7lcZtcU2XVhKy8UoYSGmsv8ku5l9YXVwyCaS
FANsfWtZWKypOVibsAip2rv2yltb90GswInCfuTvwgoRTxfojS6qudX++3bABdok
J38bGEPjmbMbwj17Ma8jKCbw7ccxRB7zh4pOlQ/UQPaJUTpuDBMwMeUNv6E6b3V2
3wlDG3FUJk0JabwK9C+MfkqIXE3djYAejkek+ecZEzIL3/AK0g2qaOEsb28jn00X
izV9hdqIHSIi4oXz+zJxKW1zUoox+0jLBloPIOiVPayE0U/fpBlZQtmitT4Pf55o
xvhOrVjBAqavAf+zXWDMei5X5wDTQZnJDF2VgOeKKEX3rbt8PjyBQn1tgO+tt3w4
dTCti1ZLxXeSnzcQwa/2FZtmZqubugupgkhJhhf7o+MwzXejDQVbpVdkTWqIS9su
mCd75735zdeQ/bKaUfccfBYnX05GrOAKC1M1S8L3mulSUrfOMIclldRrVuDvKyLo
VmluhO8gM//BlDe866H1RIcnk2XYwIhI6uX18+BibMYmHv8Fsk4v7HxyjwbOJ9j3
6sAzD/3V4aGTOfNqZN+ZY6muS6VKU9q950LZYxAzD4opb3VHt5sbwHA/MLXpXcS/
Niz3wa6hik7ZAiLCBYjNvNaMlHNiRR2iMjYvdCbDyJuea3ktsvI/AwbdNAbhGI1a
8G0akK6VB7xunn0z9Qb2VZo4AQ2fjkiCn5ZEQOzJKx8EZlX12RTv6N/kiUojn+OM
MYWuGbKBz9IdokpA/kxpGn3Ogtfx48BB+x3trL3FiPzJme8BOMn7SrH86kw83DPb
9hKeKKswoeNhIcBkVjyFVspcsw2VRTZFZmZruxOMTr2E+3EOYrr3yHZN41BL08Vn
pO/Niomyp5QeQwQRNqbSlaTRCh4nQWdz7kW+XFdmQA6ZAFU/emWPk6fxXO9SuFSh
OkzhcwzcaI4r02xgyNtxHorVJrns04Kg8oKWLIWiGukekbS+8EyjA7CsyYXZsdVD
R+/DSnwq/TEArFfY0qXP+K6CQJWacu82v2zxfvBj7gWLnhPb0MYZDqWkmhOAucmM
8v9nmRUQ6ghtxfdhVUQujfLIC4KW2XTB3Va1KxX5NYkcXq8RyLBm0pzJgCFYe3SN
tayML/i9GEVY9RBskfsLeRhSPeIHFfrZSgzFQISAru5uU30Ys3Ndt7EHI4ElC5Jn
VLBkHsgLiz14du9VdOXpY4Tu+k96UCYbdOKPqGyd9BcHqGyerDqUNQ+azJapfVF0
AxVYMuL1XILcoZB/QxyivpJITLLZYrZpGmLm98JUuKEm0YNv20lJGneZcc19oHgI
DSsbk/MkHnqmuVBV6KNhtSgq/feyhlV3NugvwlrksyCCpyH5+l/JFHcCJdx/paDD
JklYmEwOTsVshPAhEQzfkbNoazXHEfuRIh2sSTpUcVcRHtGDhyHMqkxzl/s3aB5D
pF9ca6iKTmgKBXmXWifiES/g/eCKAEPUHeiqZe6rXGCrT8P4dSntu4u7B+0oSd9Y
Sq0omVSA9NvNiGiF+fIdbkfmRacbVliyTHtFHpaaSadUaH6qi6DssPD222AN48Wm
unvKSekE6xuNR6HJ75yRrV0tYd3zeuVVAfHHOzSQ3WQP8eaAO5+30w+nZShLjWp9
MHMqJnPSNJQamfaW3nsO7y+0VHf+YM1FzHBK3QMgKIBJcGGLCtB57pVN0JrZ0dmG
sSPet0hPWXX+wQPzacN11NYf6mdCsWlgqmFY/94vWEcz5AChTwt0YzKYbud8rSSD
l6bggZENtYAzwu7/YABSRQCN8UIGhyxtN3Mxmj3tbLIpIroqoWzrIyaqLXwr10+d
1t71Cykef2T0AbR9AzQe/mNJclGi+AKRojCo6Esz4iAaLEg8nHNVwj+OTRqU2mC1
6GHViDXSZiH/KB5ehj3oo9KHrY5SsjBNyfCVU+BIhDT1kRZe4eMzS4AkE5Arn2dX
m5t700JyaURae86cn9NdjLA/colbl9kidX6v8jOIGSUgnJwawP0QIVac52/1VmJy
IuHALpUYs90VpN7jt85+ZCDRuEsQRYkZ8A3xEPoiWEytshzf4r6pyX49uqqa2Q9I
fS3hqPNay8v7deJT7DtLP9pEoRSNeV6JsbcKJ4H7jhpa1llkK11Std7c63d2k9/c
qnpC6DLTvWNWelAVZQT63ZraTFmwj93APhhbX6OU0tWqkqF3qtNEuWfZC3JxwhZl
9V6zQNhW10eljk2D0NABm2M6oflKYW/GtbJ0lXu+ukixVoghgg44JMRt3QJjw/MR
jB0a4ZBqHZucXDZYAoDJnPb2lu1uiTDbSZpc6ILEaRqQNMIYdiNfjHjMJ+3HSMuh
NG5GNEhn0im4yKLG9r7XThUOOsjA3EH06OrjBVu+qT2DP8UpnuB5nKSbZ85tL57J
3Dwk9dZmtuvlFjrGJByzkqUedsibBwEj2+rykQ8Y8rO4McArp7xad/R0LWRpJIbm
bmL5jiIVwGuxYMhkjzVNLB7eRr00Vz26Dxqxn5yi3Nxy2DzVT9IpTG+hzJHThieO
S3OxxvJ4EFe6n/xeat8Cxf8hy1D6duLZpYYPRbfXvpwrrPqd07vNDx1xgtNh1Lll
sS2rSyczjK1OBieXQ13C/ItEQyfbd/dkeXyalY5b4lLiNItJGkKOyWU8Io7wLFqD
jMY/MUCsuMXphJZrp1/OHaomqBeNiormIThHJSm+O/DHDLS/qAitmn0s5KaBRJme
TGQCFBJlB9qWUgGZ/3I17zNh6qe/HE9mdMHAlTPCYGGdRSbEFA9rHAOEDin1Zui7
z4zEV1+nzt71bfplTMe0/XveqdX6PiZszjGcbabxv/Na5Z3Q1P7I/OqvigE9hYDy
Mr0PtfMA4NY0VfT2fz2ClHdZzaynOtZ0AwqzsNGmt1/TRNXZ7f8Vs+IfuUC8utwo
YGhyViEYsyCsYR6HxTglf/+Te3JGkSeLhxmMT5CkBD5ukB4Vkoyk0rpyXXfolE+E
4syIghoCS9I8/zmaNk2rWvUQuWuvyh9T8rnNVGmjCKIZcrUFWlU/8QLLO47r3/Lg
NvlqImkWz2YrIrKlXjXtaQWa0XxD2aGM8OR7BFJAtj92RI8t20BOXDWgn0A0RwxG
dVu/PPD+BnVEVa+aWCeigoRIbn6zlPJjLEEMez95N8lckpq6WfozxuOW4I7zKgpg
bo//Y9RaGgnryMAZTM23wmbbQH7JTLHFk6g9E3M2Mg75ah2LaTyuHXxcGzvNZ3RD
4KIeIPnyNMYcXpyWNSBQkHmhYGzup1JkcYtJ+RMRcDp/adZ20ErKciTFj8ani+Eh
NbqX492NJOUXjooX0cZWmR3pq88wFZwpkowKRPKuCRDW+Pb1lpDfda/AVL8EyZ4k
TtE1/Clx+X8yqj3N3xJ6lEQ07L38RN7PBPJerh/cc3Savv7cer7PW6f9jfAbcYJD
FHBhArQu3LaYJailqKbSI81P9wxmbDjW7tIiQqVeim+QPy6RaPVfYPo46ybxiRGP
MK/QkpA0JF0B9hy8P/XK1syqzEaMOsiqC7nDyjhFghOxw5WwUMaX76BxkDyWRx2c
pV/qPYEu9BR0d5lTlBugXdwE8GzgZcbXDqVjcPcfn/VEtHzBXjRGyCn3Dl+JH+lQ
TDzxGdjFig4qEeQdEtQgpgXeFwn2rOQBDE8L7rvuG6Vpl8kZXe4a95ZCTlCqI2SZ
LcstxwYsxCwgKmeSLJ1bzQUxeLH72mJsWirdS1ADMfzepD1MkKRVVBfZfPRXum2S
3kSC9B+NQ2PYcdd1LlDZt4Kn2BENFf8wHdQrHUKg5o5Xw6+mTZa/MgamL7UXYXk8
BF0H9MCI2Mc6UZiZX4qlqIJUgD6wx5NONABhq+SS27E5H2G3au9+PMQDWXSUTjLm
7EDWIRo+wKWe1uPNDZQnUUVO/jOllsypGrYILViCwgBUTe+9ci8CmvNFSRzMuYWD
frlu99FnepSrQe/WJCdNLp77/s7gIe2x3k7MSHhW72Yqk4Y9m0MY2rRUBNn4iKow
W0Scrl/wQBWpmhjyYrdd8b+5jc4Ec0Np2sHZf3VOpWIZ6Ary80PSQIeOayhWf3gO
ACOJn6JYjgaLWZa0qW+e4/1Pv0mcYRioP8scFPH7WNFBmi4a4EQBJiXSkur8JlMv
qEpR43E4GBSsmlMnFV+klymzROq3mO24xE5+yRBPIL6/FLDe9jvHgNI/cxYRCM3J
BW4C+/s9ZMKTxNjJnhhnl4UijkZXm9ts8ZlXSRIaZ30xUT2CEj19+vJ75Vg1fzK4
m/x2u/EJ3Zkjycbw5c9PqD+1URUGU5Bil5yEpuqBcsWGXCHmTbmlc7Lcohi1sfPX
LVjpEr1QSsuh/Owhd3XaUX9sdpo8AnTbAm76BMVpH/z5pekxzgDHpufh/IEIQMEU
NDID/RRgjJM/jCmhJMojagJfRIGR7b3baTEh6FWdSAxd9PR7MeFQH51P4FySHfyp
8t7I9ACMampKFJsZ9/FapgFZcVYwU/mJn05K9qvG/lwQEwpsTl6/z9EK3nq9yfG/
tkJTd8c8ckJrjFad2nupBU07sWHTm7sp6Q2xvpxYQtRUxtND/Vl0i5rGGvsDq5V7
x5FICLjDvm3VILg+38P9yguXiSB8NfnORDN9HIPq0+IrrBYNCGufw1FPXkHS3DGU
utV0ecu0RcJwkBeYmjjbX2xtfBwZ6jS7sxjMsthesP+wSkOCCIQ6YAectEpYuJ3R
61jJ0C40t6MQbeaOUrKitgaNHU6XyHfwKQI5r2wbllD0dJ4Chb1vOj/x7f/VBKhU
Sfo1HWHU43rE6x29KdMTlpi0G1RTLu9R05V9E+y0aTw16kwfkK6fYp8JynMTRxBF
gUtYt1pTc4d4eJmmvTbNF7uBXWrmDiHwl6NrMQEEcjdYZ3yvQehyzeRNgy9YeJEY
nCiMuT0zj0MtVieD04Pq/Rn8xB/p99lP070c1nU19GQrgSvALJ1EfTt4RrVSfnxT
OFuYRURr9tPtNMEfx8JwONQYp38l6lBhK25CQtUNiGaHF4YVjPvLXo0GEY8yWg99
IPunq2WCW+Na1EaUnv0PJtT2+LK55tCUi0jko+jxxDy5xDlroMjwO7We0srGVJxJ
NdJQq8UqhVeMhEWZN7+JHictPlYwc1L7Wc2k+socbOwdF/2Ln6v/q6lt6MhpVDGD
89rx1gqfYFMSLk61kBsbP6uLNWFBEOpHrPQGXYDCxsm4wIisoo4nx+/ibqaI8nwx
O/gX4bSrtP03SvKtCqc2WHayAFEEoF9CmeczZWhFLnapFQQfrhdclq7aPD7lt2PT
bWrcSeI9u9Bd2SGEZS61a+txiDB6U2JW5lKiIQWI/G/pjne+8aPHXoT6vSXCZW6T
iuJkmdfeMBnGBNiGd79BIUim4Vc7kHTyCRD3R/3DK1bZL602KRJSDPxC7dFJPPal
srvsOww+Ex75mXR+nOaHj21ezEADi9CSNlDo/CyO/CXgaJnDGNYYsJQIPz7HQqA1
XWp0i+xN1JyTQEnEe5cjo5nbIBP9JLe1W0rHcll6/Rc19dEHyhp0FMlck9RmGxA8
YOq+ZJ9twJcuvPTBC4gF/AS6nzgWuYqEzxVf9SKFn6M5vBEUnpwTD6oLUSn99McB
MvpIzgYAyTSd2oNxjTe3O+Uurd7B0ZQIV+OMLPz1fn8s5J1qS3sgURl6OWKCEk1y
HVwPR7p6hb8epFeljT2daILCg7cTvSG9MSALnkOZPNE/MIrsdPnLvdmikTlBAmdX
4yfzp7G9O5ToTSh32w2kLFi9oo6imtmDq8NdWDKF4RcQig6BwsH7q03d+VbiAGAR
AKZPUVTahzGa7PqSknoQYKHKda87i4IHygCurzrHnySbYY9vMXInOJH+NARn4i+3
1R18JuUg+nxWFhpFm0Jz6gKM1I616dD2E+uTeHqELFcd7mxqSl7YMEOGMmDDG+CZ
/qaEP7caR59p59ySVdzwOpsNXUyYc7K3CxCuyjqF8x7argy0vJMfrwv4DJdY9bcp
hFkIVNR2q3q3XTN7myyy5eAQZSIoXVxnCp4ApspbumlKjxwGThMDOtiJrnmGwg2x
D3ca4/DQZdkvQm9z7583dDuSD0ChA/DyKjQ/16kl3croVnMBuCHyz33DPoPUHiYl
n0thWC0BP8L5ueYrHz5s2Ewa2uUHXOaOGyHXI/tWuhZ2Gd3uLRPyrBswx5qtHnwy
GKU69O3Y/2yzXr5FmYk1ny+sUniy0oT7C5P27zS/4zZHCpB3M0tURc+jDANuCnSh
Yyo45sS0oe3kyZ/LVBzziQRVKuicfFMMtDTmd5Mil/Sz0p7egfX8koH77WO9Ad9+
3xopQEAc0LG1Nlwzv5//RgDqr09VqfUMihYclxx20Rfj4u3kvSzYfLvut4HRmCwQ
tP4+rCyLSSEOJuhVo5RxpWzu/4PTYNLrvTB7hKDqPA1fN9+B/DFY/SkVmC96KaJU
FV4uciQdL4JWBsiMsUj9YJFKuKGZlAwKn5fA8TgCs6BZpzfEtXbqtLe+qHkeoN0g
zXYdhGcPIxtGw2IgZb2QjniS0/nhjQcQebf3wTy+OznZZQ0aWNVMC/fCuAHYTlpB
H4IAbN6UjOgVF7h1b6wEuOBx3H1GSdiuYoI7Bc3LmTnpHL7Hu+ywgWo41t9fYELC
CrtrGOTWNZAe0Dq0acKkh8A1iHwOWc6DxzI09FTnd8UY3LlgQQaJtOgPz9fQCaRs
2Y/xzwBgdrh8Zhtty/popl1GyCWQ2vh1mSWIsZiuD1/Y9/G7beepvYwIIO2gFsOW
9b9nLIcrO9RdxMGLRanM/FbjyXb0XqgZ5LkpfgBfjlriLta1vpHWgMHP+LGuN/aX
XCquAy0wp89kZaXw8n8v++IGMzNOkCwDahNL/yRsGccglMwqj8N6861T0M4KPr+k
6JrB9Mj2lakaO8XeE9S06VWe29LECPUxZWoQ+pUbPFekXNSGDOjd+iHqqBc+VP+g
GvGxGhrWmobkMrkfewQQTZcCiNkzwgZDs4SYB5R13g3BnCiHYK1oyESGtyBKFZVf
P1OCBZYK7CnYOfs3b4XyNU9johYeq0VB/pN5aaxK+8AGy1v80hLgAL/OGdGM0Gjm
Wj1/gpsJMwvkHsguroALZ3baRSIunKNzzPhRbXJydfUuL42+mf59GsrQ6DTLDBOh
H/j6bvjYP+lTgBo5ZMQdtZoZwN5zm5zv9Wns7sYRUbMSdWMCWWS+Kd9VOIczm7+F
DYvlat7HkO2C0/xjB5fQr9krB7GNDT+VLgBfPmGTR5YgRf0frzZ7WnCSOsw5VzoT
/JfJTv24OncDSZusL09a/F8vlBws59ZgrPrc3Xi8BGudP+kQBUcIVJBhRVAuebDD
Jw/xTGTg/gLNUnSRauBglsORSakcXXfQuZakQ7ULAIL4vfAWX1z7FH5NzDRaWRRC
LuPa+QjgeWXeHsWfc845SYmU2t62skfGqZ5MyFSv+b7frsU9L0OC4Wdpi0YXbZBH
3jxGp5Nw+/gxggHyp95zwTokdkm7ng7SThDUOjXGcxf1ewVq9ggxT+JvamIiRvRI
yUIDYkggiEQee/PLc++9Y+oYBl5FhOh3MrTpVykNgazrIaK9nQ11yG/DEADNVPL9
S9UYy0aorCugYaKZLVfwUJxmdOYvI88LLfz8U6jmqLxcKlxfnc+NyzYMbyxv5ys7
7lFNzrTyBhRyxQg7NKo+Z6Qg4xiDxRGDqSRuWB28iYggsptpDTnnOJ1JLONssE/l
TyFhue+p2KFqf7sKksFhTMVWqBaeHZUUqGqt3PHDB28TKSPz/dTGrTHJFy0v6KbA
OIMpqAss4Gfk8nnbA4a7XmqSNPEKDCebeWgOuUBJYELYvAbdXaOwcdY6iqRW+Wvh
QOETMjvmAb7dGnBOiBT4G+3nsWPWSQk+IQwt5HSL9a+7bh6T59gKGzz7ggJBxjWh
ETPaMZwfINDNuWQk9sz3EHiBSTYvbq1hBPSuD+jL1Hq/vzSecyT1PV91vE3o/CSe
IPwBbv2UKv7mFFSBJPIL6E7Y9mF8hkIfuo1FwOdEZLlDiLn0RPet0wk6wDt4scmQ
/w5NwJ947EoGkCSF8mg/jaLwlaSuGtwCw4hF5Mu/Qg9fIr65dUnL230jFUUSwiF3
vr05805bMhClPYdSw41Z32x1uhE0Qds6naBvvfZV8KIfBL/6XzkwB3sm4Ak7hxHD
h/sfNRRDGOXnZl7q14Df+E7CQVLhZrY+kA7uVxQHTBVljpizJuKCvMXn/7KQnhQa
liBPhdXFuez3lVcGBGGChpOLi2L+lAZSfJ1vBqAGKsK9UI8XEzlpRQS7iQr3y03K
Vu/UERrN9DcxSaBBGWmmMA8CahKS0/mODgg7Kp/xS46OWbQOki4fIpdwzw1HAbAR
s97BZsnX36xX1e1Mrgsg3NtFYvR+TIHsOz4b84LdBnbtSBHKRzEmuQKAtIeHQuNy
GkhQbaKjEr1HclIh2fRBdmgr72lghphhER4/OUyIo/+jybE4p6MiiSQ6U8bva2MC
/RLEn1Gf9DxFJoE9p4Ee9z00lxvEAu8UPKDJIJxuVuBYeWDrQ1zYojwtpFSVaqHT
IEjMQ+ttmCfMmDX/u4I8Am0vTYJfvBqE4zfL/RhAdWb9i5/XG05/JzAFXOZJcUPp
KumKhRJO9KF3TBbfP8D+83meFwIVN/GSfZw6LjMpoqNgYpcNei5B2G/rK9ar3QUh
O3HyGIjCwRMtdYm6d9eisxMaBNWiBN3/JyBNlaGZ8M76N79WaZeJ0V/d53wIrRDr
Xd12q1UefPdhCk2StvTCp/R8VxRt8czAZBJoVzwLzZqGgoxPOdF4C+hksZjv160I
mQPCxOYSetYakCuCqrFHcN3uY8T/X5a+5+NF272TBgc5t92O8Dy5PP5jaaFNyoLT
3atV2bfulxseQe4XqqwTP6V71YT8QAaWwGSwFz0pTLi2pB+YlpIg4VaipHrY9fXq
I1B9VHC+pBZYBOvdtHU3g84o9kjDjAN+fxRQSkJb8GAsf86y7v+NkTA9BMyjotCj
+w9A9N0k7GbLVs6VU8G2dbZOCQMA0CNmxpSKKh53fxXffEtQw1YqaDoGFwqdO2Dy
J7x5pAAT+Gov+OAVpUs28J1LMlx+REr7BgGuIKtqj3s=
`protect end_protected