`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 29664 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
YachDS4bpHRDzLXFQC4CtQKXPk3xItizVGq3FkssTW+B2Wob1t+lrTUeJNoDxNwa
chx95B/GrtvWlj1pp4dY64VkWGnyun4vEUkYECYbsmySBPxddziUCmz95BfsWaaW
VhyR8MDDemMlCbcScO+hYXw5NCH5RIRPKn6CX3AUT7fMbLiUVcMLihRrkFsd6zmc
zLcShMxLJsMj1znOTG/GZKHMtbENNvMRBnxh0+ke+9HqFF+a1Wge/Dy/ODSjM1Ap
33NvFz5vaTk6O0Drl68OHeVaaQIpdNfsY0p5UOJ0raKY09mxjCH11pATl2vJ6lCU
Xu8GV78FqmVLXQXlT6XmVp7169EiRm2le2npoCDTolOS34D31RaCSuhCs0hOL80M
280ZMzGOS8vfkCwhrgG5GH6PHNRUnkgHrYhcEmQ2QGNOgiIKtizezmK8eVPnliW/
M0tTpL+51nkfbPhC+8v9GI4qxASww/b/HH4tX0n/g0QEperuf2fGMu9QgRCZslbT
lsJE8FtN0Jcs1OFC5CDMj4cBzEkDOBT9xZP4o3QREF5gexUXq6qIex0yPnZ1NONi
K4nxpnQWCKOrVdhaFmLcW0h1pPkNLr4axtnLAtaqoVyj1JoX1nZw2DaKiqA5eDeK
KYk0PosDxAeyLJ7du0OGhLvZltcs16dAiiKW5deJlo8EeA/IlEG7UmrVNAaijVQl
ylIIFVXu2P145sodf9JcSPpbQ948ltw8E1C8W9HKQHwKlZzOpJ91rU7k4WHi6Ze3
HlbjtnHFevI0yUGPqmaEQRQgDKrStY+/2LR/KV1xrVHvRpTjjGwuGSgBLos/A66n
plqNVVC+vkIspjUsI4zeVLHzqEkFGhE/uN10WoevC2h0vT/j6bnfFf3eGay1qG1l
d0jjkt0gkf+xYLhi/RbPR+mUbwTYIWW/GQStgfPlocqmBtees04CDv5igqZ101CV
GcnPKahtdRH9UWGvadPPwt5FjoWVRYJk9BOH3G6S4yo8RSNzVby5LPCCTMRcg/5J
cvUAZAfVRuDRcMy0yr7peXgDvNTZOKtnF71c8y0HMwa4AOP5o3f2qqOs6t3Oqt88
b1HfpstwC0TL4JDCBGj/jaMbyAZjUpneyTWUHCJ169sLc6ZbbvM6xNu1OyHnIJ1p
PMKqUkGz09tnmfaqDlJ4bJbFfde6AbWvKUTP0GouPBikiCUAxJHYJkMuu4wa5m5R
r00/v3CvSRchOx6kOgiy7nGQqH9SrM6cDs3q21WL4css965h6pDm3r5ghoi8DCL+
PUNNYCT8bZIdNTcjNuJSNKnxQB0pqV2mlmvXkQ1jYbKyZFIoANmwsQH+UUuzOa6p
V6diS73r/4/AzmN+ZDPGQb0CCVz1OK6i6qiHttY4sNJtpj93UkwgcWxTYVFUgCxk
HK9zyNr00STtOVs9tnPq3AG7F9guX0gXAm+/CPvHE/5FcoP12MaRbDvIejYZqffl
RZjVbQlZHqe4zK2hf4LB61kROdpA5C1n1i2b0nN0Sggt8ewpVYfg0Z6CbBM8Nm7A
PzO5RkFPfg3Dgwr6k9LnD6Yv0HysguP1AuHH0kKbKwA2VK1f0Og5Cq/tGlqladm4
yBRPC+Kzfi0ryZrEL1sfo7raiBTZqqqMUYXbN+j74LmAOfQBtRsaezpi43jni939
XAKZDl77xbPsbyu8Q2Qi9w81+tO14jNDh3pJmmt305KfgNT2qo1OyeqTugHEx18G
k+RJmQMvwNyzzwkuHaoqSS3NVocT8twQrFczOxvn0tbqzReOPfmdHqyC7lLMl78a
c6PGRI1PWzpSBS6NjCcFV46XXiwRRxoEiTqbuL84llhf6Tlbje0tULwpml0cNV10
VGzePqz3WE0zzc7Wb2tzaI7Zm2NQQF3JjoR6G1KY16a14RU4LrtV8oqGLbni5fV/
sPmNjnUXJucMtq/O9lpJuHXnmrjwZtHfK/g67TbIpYF7LGxunORZ7LU/xqXdm5IM
cHxHHvTTxaDjdL3CcosvYU4CnozutG/9x7GhMTsTtrYL35z6Azu6A2pmnUKZBIfD
pmfvr8WK7EuFF7v9tD3gfVj61L57xJbUisSr/6cyB438f1J50lW87rnqZ9ju6i3v
0FbZGvTHj7QykF0Zn/7Hu2olbBdEvH5hWxiYrr4UBmKBBmyphQS5playRX4MB+H1
sa7EacezJGPntXNd8ZJ0EoJq70Aar2xpQfrp60v3W7Tdxch7+JOB6gLDY9fcGHli
2oGtARb0uK0Y03MWg0wPSvVGaApk+fzz90KR3OW6kqDFsT1x0zb/t8Ic4Wq0zuXb
04lu89NG+6duo9ABEWrhXVPCVP4pTx+BM4mWddS18U/67OG9nMNi+BSTXBPjKREe
wqnlTJOuaaSeCqddg4x4bXLgvhIeFm49bokKqJsGIXuHOdia89i7FcN3MHWfegYl
nqK0nPbWKWdJmpfAzwUHtyz1BcAfJx17g9rwXdruRvimBSAu0ZBBEQbkrF0fZ0fg
P196Xe6js+0k0yn7WrByzhdFxVQfhPHtiMgfEZfrMIs1J0hGbR+3kFIH1FiFYK2b
4LLsWNPcf0gE6yclyHYmZYuBZl/Af15444iKDt8XII2Mok0OY1BPjPJl5NkXcM0P
Fj/leqDoLqSZvtJshq1UqMOUQAXvX6AhKMrmic/lLzUXhTCTqlyrSmwIi4tmwpWV
kaYEI14SpeeWrtld1+qRdOGQK4NNzfDxQhK1/8aEX5XOwHk1AHjToClGImmFQF8b
EOIWydB1/+fZbo+EMfOnoNzKpXBeVfgmwb1Qt713F0d0fbXeyILHQSV0qCmWmoMA
7fZt6bYLLwAkVkIWKcGtlmfaH2DwPDi3ppn5nm1Vez8no2+aPlxY8a+WXyH6PmiE
xGFnmlc960ZkRceMP7YtDanP0xuILq9lFltJGB4UzWY5Tc4Xrk7B7lt4fO7fnELy
oEZv2W4exeQJIwlrmBVTi2sGBAwhqezjDBLB4GNDSwqAfrSBl2vhN3wCusUaLBUq
tWSO+y/+ee8OmaHDfMVLagPUjgiZTZJ8a4uMvMddSlMOpFBNyx3da2FY9CTbEf5x
HaL9Hc8gv/POJxIFugoY/JgbCUh5f/jq2Z+n3KaKvv/5PcTDSteCAk7vBbBlQQNC
ur2MXAIhxiBz38Et2ILzB+bhb+JwN8M0ZrNMIpcJj2xk9/O5ygB/0UY95mSb+AFi
HE//Uk6SnTzxeJ1TL1SdopzbKCKF8lvUEktxCmisiOErkI5k6Oa01AqEXsvLEx/G
2AlNc87v8JligMPNo5ElGwEL7ej8FoxitudompdENJrMmLh7weSzG2SEEmY3KWrF
Mo7430F8nZz/3irN3WrFlW4hWhkfrxC0fWnXDLnNORmjPz1fpdHLL7tTnRKLXowb
oj4C53nqZgiFzGpgDLINz20Zzg9PX9jpo8k3JNDmofK/2XxIjxg/029pLbyIoXkd
SWtPYhZO7BMEvhBWRZLGBdNBCo2AEXwR6qDErIZe3aAAiDqNh4AX5F1L5uaTE/6B
LqTkpxtyANV6CZEnVDNEV1pylwCjWSU3C/HLomr3M8NC3O7m209Fdi6te0sqzTFN
LWt9saaAiHwioKJ0rvfcRs+3T5AGaJQTEYmqtcFPGL6vit9seMHd7Lj0Mvel16hW
UEMDcs4wJkh3h9bfyLUsOVt/+lVppxRzA4UzLR+9xfawcMiIlv15W68AJJsW0zJK
ZCNQ3DtYbIKAmnxvuj+USoV2tvS6+ejv1E8sNMA5JoLATngB9hqb+Thc8u29hRFm
XGhwnsXoiJsE7KNdQMrWrN4woSYHEHzz2uqal0WCO6NIuOGDSVzzI6vRpaAy3NTB
3chNBdhmLaY1Nrk9iHhHx7+h6bYiFSmrWdJyFytjdamG/kz996pHReVQZNhp997e
Wwfsglx0jN9dYkFpQpzn1Yfg+tgF/Ad60TcX7hYoCZ3Oco/IUITcgXj0o3ok7xlF
VIQyoxfoxpYLXUHvmYXsXiNeGfWTrATbjViwkhKGz+ekSqXHRZZvI7GY7z8IhJIU
/jLiJ5RSvkqmRVPa3wC/I8OVwROjo33/AQI4GPTVK73rZTs8RDepeDxYhF38a4yo
2VN/ZG4P0hQ9c86+z5tFozXkTG18P6TF4Rb8b7Fqz5s5xaVW4+O3D8RcDLCY4i4Q
ZbUT2SDxh1qyxG88BpSs9XhGjn6FV0lTYUpibrsi+2KhzBXQmP1sH4Pl78GANJnH
cRa4pzb9U/+v1TiL+jA4HXY+yXfzYXhbNIBABqnEcqRccURir9Jce700CvBqDEbh
wHQXG0eXgm/kXjrUZumYduAIgmkFq8tXKDLmxet2rDj5sLnAZsxiJoEbAU9Pu1Sw
aJ1bM14xKWBF6K5SphRqisVjZXE0wX0YJLvls+r5ScwIVHMNnVg0LSCPsVSJbQIU
DrLHeyhZoNYL9oe2ZTKnv2VQ2q0OjghHtbQ/KH9Vn8Hx70LmjSe561orizHAIkVd
3PVoCdnA6CzugFm6QUUrnbEn/jPDL54FTdLEtuyKu5orhv+WMDBd8gekEQQ5x1gm
+nCNMHA0QpgnBdhkI/NDpTT1pc20lRgyefNRdz07t2jF/aGyqDEKfiNnLf2S56nm
eDRKfDLZVD7Z5K7wejD91cczTi2V6bZ7MJZo2qedkM3mu5LPeQm50vpQDO3iW1oY
JCQQZnBL2Q4bzjJmtdlM8iwMI0MPIJRC0NlULfNcPnXEQS7PILC4yPtFd0lkH/+I
SfVqTFzMTseNiClbBZAKnm+2admLqyvWapf6b2pzBwK/sC5DilG14ZND+9W9Wgul
seVN2jxtJuooi37ZbYsDLpcsVoeLI3DJk0ysrQHU5L4mBN6GcreOJy/stYrmpYKQ
mlvU8TpKJTv2GFlFgDawrhQW0PXoozu+tV1YG8/ikl4+6Datbav8HK7LrDy7CNSb
eT6BrjQuGqwf/LMN63RiTBSBmIpbYYpJ0Gmz5LXoEjTseZHTw/kyxYoCPXXehWTn
sxuBch4nY20LjNKErXTyBG8hsgJWT6KicAg0vqAjkR/OzK51Ypa6VX87OmsAGwnl
YSrnXsgDGc/rr6+XMcMPvQHGuUzukK7CO4n0KWrCrr2nvQL7mPgAppU0WDC8KK6i
VsGJi8dbva07Ctzz3inh/9aJXYrtAD3Fw/RK3uebv24yjBe2ljAWxtH7S55pgk+u
y/7DP6nuaGjgAHsVjZRa5Lgo9tF141r0Lh/j60mnupEqwEkIFvG55ORgowC2D6Gr
2hkgxkfqBojhLB0q8N1VehXV4YrFvQIq3TreBmkp900wbl5TPh0R8xudm7YAfvsI
SEIqAyLbfqzR0JY+2V4I+almNCak40iX7IywYAooQ2gWplCNMYgzp2fqevISe46i
HITj/FjzUJKCHiQjFiIidIbFd0ruvaRNSguqUhG6wbZ/WCiaWeTAqJM9J2BtLPhk
JKHL94wE/eM6qlaot0jHIXZx1j+wX5vuW9bUOcwNMDeZkSiDtuNz8wViZNmIZP++
4+8/UxpVyJUeRsStx6AozWWoIXyCth7Z6+eNtN/81FpJAv3gyD+K49lKoHnKb17B
KzX0sF59jcwc+qUUkGWtrKECpN+u8FZxiheojvmyi/dmjLcZt9aSxUbvs9IH9X9K
FBBokQzAlyeqsmvDmMxxcztUGRWr7cjgwSd48FgJHJGUtd9TB8LnVqgGI6IDY7Ut
3XTofwzeIEhKmnvN1k/kKzOOM6i1e7dbdPF8xnwHCBOoLMmpgUY2BbKW6nJgu+OP
d7w0OyxIAHVCD4hP2L2DRS2eKNVqcSk7h47e8MpCyoDqJLwj91fGOwcTYuA0WqlN
yXVuBqShDATba6ahN/cEAzjcIBhVay6jT0676Hqv1sIywTim0lGns4ZXfTo2Vrf/
ZLhUkAl9OJcL+ykr7e+ya6Xyd4ICYIcu4937/ElYwuHqhGqIK0554UevrUh9mftp
qk646X/SywafZ+p4UryTdCXowq7gmSKUV+/YguyW+PJxTuvvsugx1wPxHC1/4Co4
UMYWXVlr6ooVCAUk+Iw9XyKX9mLIW8hlaU/IEAksfdAxMDiboC0kGsC2jNhWRGAV
JYESlsl0O5o3T2MFaiN+VMVhcHSJzfoSF1nPlNEVmzPaY8ZvUChObOoHij+TRZKW
asNYqYrAqVnVFh6o7bSLSq2gYoLk7chLMF9qNx7+1nqwZWc1FAUzIBZLZE6F6Yfa
CpL6kDV+EMLdcJiBsWdFBGb/RympbGic+Qx90Aw7bjuC7YdI1ya9r3Ikaa1cwKXS
199FsZHkkeLOpRvV4/2CtDKhd8j0xG1XvUxDzTz6gcaSMKxPuJUX5sC/nTJUgx7r
jdJp/wrttWK5wetOOFhg8i5ppqyBeZ7DHtq+JYOqxYYD6u+kXLO4IjGhOhKaBH/J
59brBCQs3o9ALCnBvfKEYkICnG6Znibvwuh7KMhHU3xdKTIEDFAXufXTUjYUPzws
/7/ZoQ9liuSAGvrxeoGK6QBWa3zZxrtrK/oalcQ/HZAg+1kq3Vt6eIDfaLPjGifD
toXf1keX15pZOgq5QXOP/RhX2SdQDmDtIzdmAaUybnJwQnddUIf8MckcLjvd8fKq
4H3uSa2wPvAE+RIYPduck6863GfnocAj7TZ/GJ3sEDGZ8fJ/gDuybjDrBG0hBprH
HaM0tKrwtR1kX6EkYnLc5rswkbX7Rw4LazVBQpAI7SOHAALeSeU+w8CTfU+58RMF
PRRKmTRfUM/bIuGFt+8l4imsRd5V7J6aKJk9BQz/vr29hwnv8oDvaDEQo3vl5kWb
pE/ma4B5LdocDY7VWKmHjh8Z41E5KQ6z/VWp86OxmrOIhEhyyC6+VKD2d779SCwG
Kb1UgFy3QkdX2OuwZC7iWClOcb6jZ6KpgUsZMNtDvb/3wzWIuSNUfVYAzpOOHa6B
lHAQwbeD566a83HJgKGb5x+a5nBMnKyw5oFopS2MATG0/6u+kg9N+7LBaHpNAuVL
F6oSfTcA6J97vbpbgS2gyO2x/fqEv8TZGOofqpIAdrsYBAG9FYvYj2nhVaGrJQLj
5qAlrAu9/MNSU5rkUROBg7Vrzn2pUYSmltwXe++VvtWeT+g1Uy2pgM/wGvjtxQpk
SAWh6cRUV96nplo9x2JIGVx5UpASdEw96sXu+PUoWWmbqdBUzGb1USiYLvM4EjgW
pzKywZCyt+Ewm0zI/Zrv3Vc3DfMbRlRYheEPR9JhDR2LiwkgK3co8lSlfnqZyHvP
KFweX2AOdoW1DT/5mVd0Q55Yii3lzM/+Bx3OorSUr/varKQZ8EfbXviSmbU+O2nv
Rj/jbpA/62PWeSLCFXVRO4nmFi42aRIDaf4nAiiMX+3mxJ4WsC7+76EjbAG6shra
hVt97Ep+Uijs1Hzg75LwyO4nvv11p/ApzEE1Xjvd82pGvcU8p1//OwWzR7R7DGfn
oaOtCnC8XRYaGHfpEXNOIkPfMSxI+9XR1oqErJ40rK6XLrdZmpHD57YO0zLbSEzr
rYDtjqYnPpBeS2Bimrs9tC0TQVrglpmpltdXUJJyk72j5Om5xDJL1cg+e9sdVc9T
frcox9HxwMont/dlrhJo+VOmSSroB+08z5yZN1cDVg79r1dQWSl0X1d03KlQ9oTg
2zfr57BSmhqdHypF7Qdl7ZMLpACeV3sBxRxvRdvBQvP97KlBdRwk7D/I8NOgYVa8
qTwrQs6W8YhZOR8rOXDt56E7Wxd/GHht7L9Eoc3SNs7FuIP0VkaDd8xSFFMMX/L/
5SoHIOPMqfkljhongPqaS3QNjHEv3eO4TPNU3Hfq/GTfu9UjHM0zMraJLbZ+mFHX
+F3ijm4htVJq6w3leQ3ECXv6S4GfG8/dIpw0FdCDqs/vXCzCMP0o6LCXHLZsS9Zk
RcFsw6yHbWiiDzgPzTD4bIFo15PFcTL9k//EfeO/poOj8ULZasK+bJvlhOROTQ2X
hVW1CcNzDTzicWXYOX4/9lVkoFeg04J+Jv/sKlRYI7dZ5QXG/CntTTRLftIkxVQA
VfLM/5yZlLDou2m5+/EXw+5pX6+53fhjxWw9zNvuruxo8ZFARpAv0CSbA4DSkrxv
EtidOaYfyNc/PCeDUfw+WR9Hehc8zn1Iit+4w5yjKhWEaSc1L30eeroFapOaEnGZ
FZVrsGDA94/0gMCbeGjmJpSbTZdX7gQ8rpMQAwj7ubq6F1YZCrMUsO+LJ90JxzTo
oQMTWiS2r2xQFQsntSQ+MtoMB+7nJMT7iiHfHXiwtMICqodkdzGfTZNfz0pxnQqO
HjdTJE5eZiYvx0n+sBu3E2RL4HRFgBFQxIQtc3kdmCmgl/2/BeOm9/I3ahcZ+5+U
RLCrrHAvMAGbqpo5pswgpfMO+716MB5mLz7prN7oW/p+glIQZXwifOxtf2o4VPHG
euHzNFtfQW8PUal6uCArcgn4kRdy4ytgg3ne63q8h6HONyRfdpx9TME7Rvqn0fsw
ZN4xRuAVn9zUixmhN/Vw66Y/+i8QJ232EIuw8lWiU7/UHUcqyAzjc4MGcaGuuVPI
Q90jXBPqe6IE97k6jXBmmnFKzSdhVqxsn3Do1wL8KGuc0mKcBC+mQMomRiy82Iba
Z5j5DS0r3HRRFQb4BsI7LmxXPCorGxFbWVNX4sht86fygNy4eF2tmj8H1c/UbwlJ
3C4bnxaeY60XdeB0WC3/e71Wp59lXqCRvXLmNsDQ+V2OnyI2ElGz08mJYdXqmN9D
09A1GD/vQ3bE9W1JWMLxTDVoUO1vPoREKorWBRje4kC632oizqDAlLGtuucROTvG
HOfR5WuT6HknuN4RrR3ldppr0UxTxe0Z9cU8azMkINAA9F6+99V2XnWhqo0n3ZzS
ZuEn/v+ywaApwviHVEtBylTIYqi6+crD5y3LxbmrdH8GuJuxZSPu4VTuAudTEURk
0XTErhmPfDkqG1e94nlcDbhiPfXej5zWsF2wc5CfvMiNRyEDeWTZAJ4w0zcOqwXI
9xsNPO3hZojT17WVgrMrOLNAupDUo+InRf0wk14gjg3m1nJ0CMzer/rJLFB08c/W
3q6RpVX1tmkYJyCIhLlx/Q9b0inneNU8EnYKCUHe6wDwCAGt48xrxRFRIiuq6sYM
5X3g+hSlL31hNY3W+X8zRyHNgbd0cPB2xzAS/AzlSP1GNbiaDTau1FEJmG7tKyy1
pktgnRIqZ1w/DWWuEZvuMJbJmhkNUITa7fHMzR6S+nk8blnevK/PbmM2XgNRP3gu
mnm3uA6syA9zIdzsYVTXETRTUkWA3o0fnjtLiPvtCPzqwUqNC8R1GAc8iWZ+SXfJ
LlEmunqmz7oVGKKpCo/YCTkFuRxrn9cPtdk2pHOUaTbHDKcUlmX20tgARPmwTbPU
o83LBf4GPyOWRwR1+gVZ1P1V35KzRjFltm7b5NRHpAZD5p16s6oixNelH9tm3jKQ
R5pq+VwvkIZRq4Q1Y/49RoCx9P4btSEfEE2QGsSCNru3wKjOidRSpvbfV88OVNRY
G0eXVMQP5cUA+tmbgO8fPuwjGdAGyugZgDe0VMkMD7kFLzBwki20OfwrblnOfpGQ
jolQZxL0LJJE3F8wre27m0Sp9vKkEjY5TrSIucuAeaAF4AnJcX7FvH+5qRAt9bKV
m6NkelDLJ4nu0QCzbLvEGv6nXdPKq0pRh9UCgElpAE5wI+lpeI+v1Igr5T82cSnM
iieFhlbjLRLcOIU3PnrL6/FjQHQqZfRWaooMKFhZ2xKNgKvbJ0Uiu0v9eTnB0OsG
7PJ4QJ+w6askCbjIDac4vF46DHC30GBxNeVv/ueq3d5dKAG/Y/v3i8dvUdVyNbWi
nUcXdKOTmzUDnDmjRGquN+yUjyCYCJNCgt38gdipkv6beLCCYv2FhBZ+p+HGDkSN
qfypG4CdncN2GB+yO6RQtct0+hSDZgr8RLczj7Xl6YIfosn1D5oT82j0YFw2Gk1y
y0GG2Pfb4ki8yEcNjAI6LbORHngIRANBg5ZM5gwZsasjgg+VsxY7QY4Uo5DtpSW0
M8G8nQmj7QQQv3qMK5FIdbs19CAhrA9sbK9TxFbBO7N8JDyD8Mbc4v8FIvx5kNtW
JnmVQU1h9+w8bOaSf5jqLoxhBqtZGICJ/uVKnkiKHgu1js4aXByHRY0TS63nJ6cu
wM5E0oHj0NaGaOCmjI+e3PDZ69VbgdjgmLeJgVBT+ICDS4fcyWYVe/Z6dzk/nh9N
xqFbvjei7g6tnEs+DHrM2HlJ2iPFaSPes2mek4N26fQbf5zXl+SJdtxX4qEidsOO
CnAbbbBmrkfK7AoTWGMPW/3A/fF9VXIZD98ktDUKdc4xN9QpSzlJI4p5Ptk39CRn
BzCPsX96kaaOoMH/jyQirmjuu52sa/4JO0NPZVcAFgxv1rgITSvRLW7+mbvXDvBP
Hc5uA2u3SZtMMlKvaUY0/3fexOewZMlhN/694nNSKQXtNIN8whxcsLGDfvYBQ/fA
3hjKMnw0TpH++E07jDS/1YcfHzxnDahezHGrtWg2cMVWCzlZsqyXvUaBpCFxcncc
xLc3YrgIYKbt0Wt3I5YVyGl95lZgXmU8HwnocFPqlyxOShcUKN/iIcPmMiCcTcNf
4AY1vKrpiXf8q1t2jEcP8WInDvkcy/2EAi1XZjJr9MEqrrFu4cmbBFqEIdbppIwk
uIHYQ9c6D1Ycu6mDfIZ++EDRZfepHj0VV7UzpMMRLB46cCYHBSr5V1Kob1ZFt7FN
lMt14WLX1OjG1rRxlvx4Ap5l9Z0RaK/Q7+J7/WrPlQGVUOZW2cjSyUcUYqCabGrh
vPjebJDlhgSTCTB2pVoFI78ciH/agowZVG3ZM3pFROfNSTZFQWD1pDbaztv/FVZl
VAfXIWL7zLbJR4UYRy1P2Xc2IylPnfU9DT6L0WKqW1w11brCYA4vFXqp9sV+k1aO
VMll/4Zc/cYvDRHluPMkMALFuwjcxMkShRYq9Sfi3zJO3Lsffrjhw4eUWtDi+kzq
v9w06Mwm00UaWToI+fcCHQcuGIcXTWxgml5Xr1FpSdf3WxonQR6+1uqyMX+dI48c
b23p6DKsSzoSvEd1e8VRRmf7eXIwt7rBMwVVk8Qc3yheVPuLBWT3eA4aOc5yg34Q
0+ZQ5yR/rU11oIV0arMf3BgUq1cVrXf7UoCgZcSwDGk5m9jxCQQEjuOVgi2DQb5A
QDIz17B5GIRx17msViHdTycBJeRmT2ZK2TerVSICLIh8LNMqgA5kit8BhMvBmvPP
V1vSsNqW9Se2VZdeqr/DGR7uI1sgrqs9KPCBeDbCux1ZaUtA8f1JwD9D9dOif8SX
UYv14Ns4G+QYbIXAs8qrMRvZNtDw/HozLUaXumswbbo6iOaNWq/J4e+mBe6odTqu
NLpb0SM7fPK7lnHQDzlwoCZEZ4vCRFZMUHpfUl4R3zFva4Hdzvy0bgMItGtk0O6F
x0pLClRzpAE6yIRQ/f2cbSeWgX07jsU+56EOFN9QF7xxAwc8IPkFgp3/LuFVxQ4s
ueNp3SawF78H9YYif03A9+H1QlP+FqXDRnR3rD1S48qhYgq9nree86T82hUzTCnd
WCH4nUK/VI9Js1nV7Z4GLA6aAXnl38ZZfZ+wVGTkXV07H1srd9AxR2lYoDEc5Fo3
sBduan4hQYuDojmn5qMyvPYMHfyvmK+tuQOxyGbHK7Sj4iOwYh1rrHlN6tXsX4bj
zR+WOl8BIa8bOt2x1NFqfr9w0ssNt23TZaBpxce8Zk/cXGklQ1MT3U225XmRMqe6
P6rtHCJiXW5csitWtpMq3OpsoCuOgb0ziexXz+VlxrIa/8VVoEN186BGbE7YYsnp
l6JCzqrvnQZI33sVEEeZcBmiNz4JxSqIkexWhR0mfTGm4Z4vfFN8FowMHjZ4OFn8
QKh8gjPuw4ZIHqhNV4dSYM/Rd34WOaZOKrxPMUwtGLXlYkkxRn0T2Rq17CHUV//s
9dNV7eK3Gd3icBGDYmDl+ZEg1OJls7VxB5234vEd5+dMy9VZ9z8rIG/j+NWPg7tr
cJzZ2QOaFSOH6H0KH5BKxlakTLIo3ohCfYWLphlJLPigyvCl+lt1oNiwDA/kK76R
yI7sOlSaY162/ZzvdE32pG1O30rQq/VUrA7YQjKsxRHKG9AAmT7DFxxvctbyAKcc
TEeFvrmHVcuyZR975hL6TRfQmFJQAsTY1tKgrSYMCbw+mQGo17+ZVxqeNfOBT6fk
FV4Vtp/hkzE5rtI/fnoi3qiLmVhP4vROI9K507Lxa1t3Ttehwr/vUQzaeQvUXepF
ND0bh2ozmuAwk6PXdYllvKTJsfy4PdeZ2LMXslUteKtUpkN90kvDZv3kh+BsOX99
1it6OLXClqFXvThCVwIsOPoyvnmmklHlL8op53OhgUyGSMfYIQDAno32CvYMtrrt
Swo0pWouHNhQ1Nsc4fQnv/z0/hBc4dwJNwtsxx9dKOwIkNWHmoSPUuJqznvTFALU
iYwrS+gHr1M2sas7Wenmy+/YmIRoWjjMjjAM6uFULFNxmO6PSFmBzmjEfXYQDzGb
c479fPWZKR7fuwHJA6R8utnT5onkIUETXYYTWIrErYK6ggZoy0jCNga8ROQfpvab
4i++dU4lbllMErt9c5rQg+WZvQcrOS6d22B6msKMIvfzcvGewAchncfKRyFDx3lE
WRE6brqObOOpama0nxhRai6mITlfRSfYi1HgAZrDFetFkl5gP1z3n12o3vbRTbSx
pzN28at6jkRA++JIMvaVJeSF4vr7gXD1tZYR2xRXt/7KKRyjakpQxp+Bou5YFIsw
rtlAIoafHwfPypixKYmn5GhxniLoK6JkfZxcC925lHjaVVyBLjP4icJwTqkDzEGr
AvDYGSsd5/i8IerhWfGEE0c0upBwIxh5d+P7dAFIEL+2sHxpgBORqzbLKTMa+LXY
EBrn0b/FhahkdaMDgACb+UPWtDvAU12fciIE1z9azAwalzCpQtpZyOFXAt86TNsR
qn991CWUyAccLtnk9ixTFQitpbyWnfL32b4HcFXtoTaVzdn12L46dz1WGevd9RVM
Fy8Ss4fBdi875SmFZSdVZGTeoXEp4D1+KCFg9SuKN3BU0oDdxyrighuU7sJNP+4+
U9kxajkyDeujZ3XgqB6bd2iV7usnY1RKsSL9dZTF/k9mcITu3HVvHNX7eYiQxNlP
eymtoevPbPqT1Q9NGpA6IJzne/pZlGwdqOmWqasGIp0gwRIBIQBxXpjUYDL0bMcF
b6Mpt8/N7PnWxR5RBu2PbuFCBZDnBHx0ZMzXOaO1hOQhXqg5AZifXA/HPLrniTie
9jN1C7UgM1xFWEQ6J3cjfiqAeWvok7GXOzM7X3Lg3hCpP7+5DNkxu9mBgTscJS85
jvN2TDk0RpxUWuwEWpIiDRs8w7Fe8DG+0wRrsbYc6ZlvV9T7XpwkRjNQz38zGSxl
qqn2tj3t5pkSxQqH5Q/Y4EkDvsArtYfaEEVwZWHUU0wBXlPBXVPgdI2N+jjm5KVB
eerfdAqxMoo1Go+sLhQ3wS+FzbkJHp5MaUlnYjcrWheSoeNzkqFT4YSQBnTL8I5D
OxqWXbRf/CaM1mV/WIPCmkgMptVWJTagELBydIp4v19/VVQkMWPj7w8CSVriWRqC
pWiniq9seLf+/f0FC4Sxri8PZavRF+TOSFkHAddiUUxH0t4tsq3Vc7CPF0tL4Vg5
P8oXzHE1D7F135oALHOH2QfXxbJSUYos/mQ7a7wLBnRvpwH/ytFynnkklrW5gQh7
e/cKzCtgYIgv6IB1GZBZVKEKI8ypcejHPhirj1RhtfbmgQmMs1D+tJkil8Xvvl1r
L0lss9hQ4CuML6qOXDR7OLhBO+BWh4pxQvIvMIWk0RcrqP7QwW0o4LkTaF9vaYPr
oYCgxQXkXo1hcUQqo9Ti4HarwwxXIrPLn1vR52Iq4qOGWEN8rEoUPSA/TervXnE+
hV3fToVu4wnzQXLtZYe3VD8mcY9+ITPwQ22uxGH3ohYQcdxqNsXG7IT+F1sUGck7
dDwi1n1xLh+r3JJUwfZhcaSCbVZ6eAkIl1xSfHzHhCyqcFwE4JMv9iD83xxhDIH9
cmPLy0EpUJqfpE4HeNroOPnrlJRlvybVQts4Wa1lqqZWCdVo0IuPiSBY9HR9YSlm
By5m27hgtvfpIvD9iEWVMMuwdaYOK6OVSZKbLt2eER+wZj8I/02xGmy9tF0A/kqu
d097YvEMXevZQtGd7uq6jVrD1HqSVgVrnA5iBCGVrvQPZz4zS4bMpwWqAW0Moyw0
3wYMdj5FHRVBJl/IBfFMwVPY+Vw/fWqKf/tR2SUO6eFrXvKMTxESC618BT8LNKO7
XsRiVDLf5Kq2QRlVfuGtBd9h0PS+evoFTmQSDJbnHWuyJNGaZT6BtfO27ukvisT7
Mf4DOCkIuw4zYEgRyeSuCFMOxwtZczufOLIR0tyTLxJeTFDpo4LsDuECWTyMTq4d
KqJ57Ye1GOx4+IDCRIigrEHCwuPFrKiJa3nxILhOCD/f6dOTbTJMgNw13HDT5/qq
I7wiHeVq3JT2X/l2Tfh5GN8TwGDK6fAWhVVBtI7V5x/b0/Sj4uERyhf+ehp8Uu+2
YHxxvB4JhojWvIKdo1SiQZ6nsiHufcr6EqJ+nUMNcB7RcG9/0Pdsv5gYNch8IrYx
O/xcWiIJ72JIR7fYpk/gFCPRxU3oNrG8HGMClHLdPDGc0pXdn7eRCNtGBbphIpR3
G1ReTngoREaBSlNU/+jsUPCHhasYGLQqFmPNLrUbQnjDRpaUYAAumTB0rxistyh7
PPyc9/fKGG6Q7dfO59b+UT33t/AlOsp15K+suMbyHzoPqHOKblFx9qlKYh1hbzFY
rd5H1E1eOgxTXYg6ly/9UFhY9DPS2pNh4a5OVzePD7HxHKn5//LMm62G7hyU0wxe
6og1sj+USWyNsca3eAkC3YqPDme5UF2AV/vo2QEaO/bKFV+XxDMLOVX46k48V67w
ORGTCueTwrJGaxtdT3bz3HcVDMxToRLfmaPD7iPiCTKaDj9CsKvNNb0GK4p7gCZC
KiVC2dKmh+m/psinfcPpCHpgnqHxJH0RhR6x/P3NEm6MMLYaVypZY/ntpoXpjspo
AiWfqBj5N1DkpXWkaLfz0FRhRtlc0rr3amWjB8VML+sunFxWhcj/4Bh1eUuCZ0tT
AKbcaMplvrXyneAkfvZkwJTEHvrYoGXcZiBAiq6jD+jy+VaWwrWP7RbKEcUhdEz5
7SL+Rhi+SdIkAqsnybvNfETs9wQpET02WtLCikJf436usAl1KZ9daC333+SEfLm8
UPQprpkthbspCiaNf+1tMDcuBkT+LC+/rlooIfuHhAop/bUoRLx4SuWViRwJD4uZ
PLZXgN3DkyMHC2hYlL5yNx674YBZPbiRzdABi/v+8cvtOqLnRoeT+k5YD5yx7nyM
J3fgtfMAhv0PuuVvZAPEzEF8s59uqM6yIbzVue3lf0RVyEZD/DLcLOa1Qqlt41YI
5rCdFukiKj9K6M+gnOvaOk6jHg71XRFwzhHuJodU8JJyaBwuzrAr+2RTu6oqF/U4
UGnSD+Aj2ZBMiJbWl/FZ0CTR4iKgZxRAv7LpO3YOqR27at4IX7tc9H75OPspJO3I
NC5wT/QrMmaRjwacXSSUIS1288ZufkPaEvCROMjxkWMdpfyaH2yApl7/GIf8+xID
7EY1cD6/WnW/MhCmb9nT+OakAUzFBwHRNGX0n6QugqXSgDM9QBlFzqfWkK8ll3zZ
YXuTPtn6Ld/VL8iRWSeOlPGj6+oDarPKUYDAsiN3QgboSjxmGLjgic22TMQuDNAL
zWq3bzimwqAA3exDXLoQ6HAdEZG8MJN9w6+xDJbQA52Rq3p7P7CveZjN81FQMSvS
wiFLS5EMEIRe3y8TiJMNPcAOv9yroBzTOf9wwH3S7QQ0GlSam6+iyQ032Mm/xRZo
FGqjBP+BOhvhnv2OwC+Iv4IQINtyFN7sgnJ1fBWJepsKr33z3OTCZCz/uOv4gVsv
hUZphHGruNUodN5fBWhuzcLJXXts90cO4dp6xOiVDrlrIfIhZ8Y4xhHpGAoVsohC
pdmtEUx3HErQ8NhUzwYIvQsGZo4a28JtcQiffE2QgtZj5g7B59vt599ac8XNhQ8C
IrdDnmuXSyK/bE2CIV+xkxtQdzor/NUTeoz8Wzmx+8FHq1HqT0rlusfyr1TPSpIK
pNZrN1Gov77eSSAG9a3qzxhxtkDvtB1TqEkMPoQHEd30m4Jk1DElWXJ+cdqiAKmD
pBz/zPAitHBYResU/mfZ5NyLz2x49BN/ciJoLHeXTdTZFryT7HNqB3avCZunGlsI
eHCDoEF70Gfyt2DCXjWaZMyCnKIARImzunNnE911E2GT9tThR7W5L3fSKT/FgZle
7lYTHlNxa9uZJLojDOV3/A/XpbKH8ZoMfW2g5g5YvW6XDy/lmcA2WiYHPdP3vDBU
AO/OAUkgR3MInop0DOqpJuNiqIQu9Kfml+pJ6XjnwEc4tKuw1ilLtYy4ePtmsQtM
wa93bzYWccNikkeknwM2a/ZbxSNDEDN8yFNACeMLuRE7tlasCEzrqSok4YafT1hp
G3Y1cbXp8EhbH9B/9CAYcJprj65pFvZP6GzibMLx65998XhHCflxTyZQsA59LljD
ub2DeMvNQLhj6s2b0+WAAqBFvH2lO6uben41Nm36ZDAzY8dWQHx6V5zTPOfTJa5K
VYDH9vJ+fJcbbjmM6KaXbM7VH4a0EptUUh7/ie9+gPabco1YZ9tvpIxeY//SiqH+
ysdFhGmObKnPFwQZJno+RNk0AVxorYzixbSIZOK6380rGTMAL7LHSQTUK/qyLCHM
KauTTfrd+ida3El/K1ifgYt09yqapllGckw03UOtXzxcXfVjx59OMw+IVQg3FnOW
smz5HqUo82rwSEFMRN3qFRpzCKbBIfwZz638HRLadomZdo6zkOd8qIgVwmKVirnS
yG0T+SBKEVZx/tunfA7zw4+VV/hUQNccTsNjBlmYXcJXY6+Alt6LMRA9Hn1rPHqw
vcZIpbrIF2C9nTtafx8OEMrMTB6boTF8jYCgsusQOOjyNzyjdJJSDA2NfLfJj85q
L2stbaWXO0VKT9TgCt6oJBKn5NZqMAotsQwUXaxsxXCMi52ZZkMoIBFwMW0GIRGp
HHreM7IeyyDWTAD9n9k+zcMcIWOV6Ck9RUK19GbhYGJ5jmw6Yj5EIw/TnylLBGLq
raPdBq8o2ATvlWCgMqSZJuyf/D996mEEnoKfzUShwCjcgi3F7+UhjfYT3UxUgiQ2
TbRChm7z2bPeghnLDOBdactiW/A7Vf/VmYDeHj7K0PfmdhhJcWuR9acGprGGfUP3
kuTMAYaL9HUxNCbkcXhEaQLC0gY7DfK2UBi1NV0jdGJBPzzTrQwSyVxYmqkV32nL
daIUWpKS97y8Pre5AhG3a9s2klASdWmbxkcbJTehzNWaMa4h+YrmUrrhA4OLGaKc
NtHPKNtYDcrYKK36Dx9BL+KW+ijgrOMjRt46exlry6W3QjBpCWw2+BZem3+GwZWo
8//Q36JMiIWSEuva3AzGFaVbn4seGrNmLns+5ona5oMMeap8/c38CPJpEYsT1DIy
P5/25jtM7wJcwtDEJXAy0NRty0zmfiZ4hkMiLbZ7MgPAefcDQyzPidWeuRaQcIoA
J2PfYTAfc6oiFqlsBX4t0X/7ync0fyTDsxFUXxHO/Xgf2n4RXD8DegzqaDc6gtBp
NcJBCaViJR0s7hnz9YG4AtmJO4yEmryaZ1SASdGaMtkVt069qzyalW3ysx48obLe
XT3nh4JpPP3cWzwtc8iLvXKUYD6B5hEU8PKvD71BG+SExg8HbMqLrTjrE68s+p17
aeNc6js1lbS4vlYX7+WuK900yQML+IXYFMf0nvRVWbEsfd1qVqvmscBxjZzUtnPI
djwl5jgAFSC6yAp7YjgrdGVXL+zPQnVk054ChdXpioukS5dNxbyPF3rmPf9rWh/c
VJi/9xfdd5B8qCwlGYju6etSwI7ImZgv+pvPu16VVRmXThocpJzNAggTE2Vhq08Y
+soUeDCH6OvGjjWPxhVRPQbo/+iHLyYohXBj6tXYLjpb1uPDqw76A9wekHozpb7Q
LQw18pKV8XHr73jRJhDsqByYjUjVFrJu/eCvjVcDr/frxqUtu8KkPEXwuZG9DYwH
aBGROvhCjhcDOit5hOI7abREWJCzek4YehuuzSUiY9iQUgdDTZ3sY7GOyissEjpP
52MN7jvmOHTBGw5VlN1gGwST6mckaOSWXyLoliPZhY7Od8M1ZSqyUOWEAis0MU8i
WcUQlc1A4pRguavtfnhMEhXWk/RTHQhT5685WbdEx1OPEcR0HIaa2h8UpgGitVS8
6hUSJyicq3KzpRj63hh0lIJwAiHswHxpjuaBJlQhS6pOf/6KaHPvJpZKgr+6Fw6Y
B66Cf+8GcG67BtKegVyKf/7LQqpqHcUTpLb+J0dfKrw6A2t5EEwnRzYW10gkAHn4
6Vxkfc52dSEn7LUQtrpjVrGtRCylyIelTi7IvZ1sSA2FuZJZCDhTf8XqBGzxHrVw
Ebk2/PUAbGGWKYH8XCBJjrZK6FKVfV8aEd51j8hd+fctv9EcSfVMOs8Gu17mRdSI
ZjiKOZNqreJ49Ig4d7Rt2YxROOlpSYKP4RrK+x1kl7PNvhIUiiDAfsaMl/ipEcI0
laBJLeXmvNZxZ1RXZxUQFHQHHnetthaGQ9oXTHu3I5PPr1hE/waPYGZEtYwcUqeJ
XyTEooPfehpvT1KzuIV6TiuW0RsvW5IiZ48uMwcphACfOqaZoLszFM4aVAL70e58
ctNxVvsSTrx53j+2+jwbswhu7ExadyNGME6+7sM+caZm6MPDSknL4oWK8zN8u2C5
LDSstCKqr4BDgh8PZYNE/YzpF4J1RwBSj5J+mkxwpL7bHEvbE8cT0mmyH1lGd4Us
Ijfp2ZCTks7TZnHFPyVb2qyZ+Cc67FbsjZ55h8PekyBXcZtzPJuotOECYw31aV+w
7EP0BGqFqCJ4lSmdbxDS7M5FgMm9Tu6AotIuCFo9C+i2jT3/oSAh/jzgwViBdQAB
7FBRrXEyrjwEUp5Q4JufLLj8v1//Fr0p+Qgq5syuFY4h481mbjo+5tbDwU1bsTRk
9XSZYwuErI1OyVZ4Eb70KsCW+hU7KlNVeYsYOIem8Ahbw8SRx2lkGvCpFBPk2+Qs
eh9Qsj5oAF07+VQjYl68lpcLJhkC7SB7dq0jnOQ0/6SWKQpeOL1WlsYG9Vz4WpQ9
sxciGGsmJUGpTJhMXV9gkQ84s3K5MdMhLeldRmX+1wfqCZOBJS9/Oo6tRDtj7Ofz
4rZOAir49SZ4k9J4aJFvxRk3z1ZPiKVclRmNXazoBi1UOBagBYilaCrRR6WgapDv
ep8SJssfHEVqXB9mn0SXBTBV7+AsxITCKg8GfOwsGesl3ncC5G9+JFefi9ISBVHV
KKbLVaRPU0QhoEaJXbgMdQU7k+LbPebM4Zb9dJRUd26DYzgNPRnS/+Eg8STBTMqe
KW3/xTjx/OVcSAkLu3UXd8JAhifwaNuGbO1nhIeXzAELFUPbjma3MFibjmEJ32x2
VXwuHAlhfifylB4taM8pMxmLzNTwKHGZxMKuyFClRj3/c+MtUL2OVJP3R4G8V7Xd
6uNBt1pZHnTc3JM2wsXdNn2SO2LvaOo/+sgDjNak7H2+CrLte60s3uAlfmFW4Fa5
e1sRveax9jGLQpoxk2E6JcTG3c2y0UychCsKIH/JYgKFWr9FuMmXLEoZ4Y3oGFeD
50KUkakw5bBnsuxvPaxFffxXIs0JtscEfeyrBzcUiK2pVjXpgaW8EO6Ud9AbYnPh
FWLFHFJjQEIbTL6poK9Ypl2DP5CO02AHVMpntIy/YtyshZ7VBJUs8OIWnF5n6kpE
medw/xCuEBdfVfKcJLXHgRErAjvLLKRnbZ0/bqsoLQfHXz4VB9HQoGPYC5BelBX7
s2c0wX6D/tByGTZPZMvX0TAyPgMoCWWfe4IXhS9UQwjLBoOWi/zEMbLbcQReaepB
76wd7QLiIFC/O28tkOBF/8lsV1Ss3ovnHIJqb1SQtXPCsciaUE8qIejFFAZrCEoN
FK1SekoHtzkzyivZTjRo6d7btoVW8HbvZwrLq582QbkClxBxIrrx8I8AnBlpQ/rY
vHHM1Z3IPfeGqbt32/wBZicYhZmPRdQFyyxv5K1A38RxL32abdmUrEvo7XdLy/cw
OlTjV3putwZ4WGXaaDbJeS8BkNH7o4Bi+gF4mUwRNDyPHmbNzKISJ2PK2YpZZyb0
S2gwCMZqy7xgp4MQdzcnLTdZO4M9+RiHzaou4BNAkrUfa8kMdgiKDGn9DSn4jwVu
SvtVFLTEPsVomjk1i87H8nEYYu6krkEdQczGQckkcI8dRsWTqX6AWGhycLEWKlsS
xRpEwrHiW88KEqOhM4SrwqiU3HqwmjzVj57jbmAEiAxe8zBp6j1TSnsrNbYySoh5
55T4Qb/5SLbYdNkKbTiYl4q7ZkNlhmaSRiih34+HiS50zJuNQXs+J0gWGtrUybi6
rFhgLbR9dtLBtryfZdqXvE6veblsNEOuInqu0BvnDqOZrCxlBOHJKkMpwpovMZq7
M0j9Ua7kNahma+hN+4M87s9uaGDKc/0ar6rHZ3O8kxgMDYJrND8rZSiy6kKzDwOD
W0DEzXJ7fPOdNgCfHsYsHGg1Z9tVwGHAIAhLhyF0KqRWH9lnvObb1YkgCn/Zwf0/
9KZGMKm4bi1E9QfrG/nCx3tfKw04U5DpVXBP07+ZpyUGSzRWHt6+EW1GeyLqLtD2
zjNAXgeKmp8LVlkcVKtODiUoO1Tgg3UyAERUNaUCqWNtACGDGtiAcAWdTTsZLoSZ
bGSnWv7+oLP+rs0CUVJZVcv7IiwvQntOd68ddH22GAKHng5kTTP1vqlNZ/ppnWnJ
0vOhKwknXJSUkVXULlwDzR+hkE1kRVuS5UxHghL1aYzvQFU0fuqrH3ZaJtxsWpAB
V6cUkyzhSQJpt72eMs7wGkf8KhDbdRdjB+XF1kxtw/1Bt00j7r/idKYDwcqDofbE
1JOcJPvphkFxoRQD6C2vjWzC16tqdR53/n5zX0Mm8grS0j8+Mste5BObphvkDyuC
T28LZo+WooK3vY7e8sZLmcJcbrLoDFaS3hF+yYrXCBJPbxsEScOQJVCsUs+V1b+P
nw0obA4EwRgERUkk/1IqJDqTnfZNT0NDPoKVMt3gzDZTFpLPRqto6EQrdicuaE85
ePB4n5Cl0L/89eL4IxGjpOMaZNendvNMSLttrLe6iEQ6Tk/jVsL3wGp+gQUBwl8y
+cb7t4IJMZf+f3/oXwx6SFdCqAPXjK3c/x9q7D7Kcl7RfpKvFfH+kqcClmsLli6K
TZs1qzbUywQfIajVvGitt/+2C5T01VPY+3q7Vs2pdvzURUYuisk8g8Oh3VmOhX5G
s5WNXnSQcmUQmcS4oMNaEq5uU+2AkbNbE2KaAciLgex6CIGd0QEGIbr+MOaSCHe0
K2yulEq8AToaBnmOepGS6RMV45KtkL5GKrVE9iQXCVwM82eRDVS34QDuA3SFgVSK
/2ZI+iRXzIUkX4UB5KcffKhuB1Iskxy13hQy40mTYXzFyFpYteDS3AoPHAfyk5FK
vKlJ2/V0PEWKeYny0Ga4f7T3ju8PzZ+xAbpnlGdPAuGPanrFoiAh9abdIeovEC3g
0ZXVyMewEkdcgRSyTmJoiwadoOGpvFDMPDLeMAtH8HrsaO3RZbJyrSi355nyCqUJ
QbiAfeuNhC9g+lh73p9cloOEAHarRljH+Z3/bV9jzRJpWFPLeJezlIuv0lIDnI//
Dkgp+LaWzp/5HDfDpkR/MZfhIyOwWS4Gh3jLmkROSfXzKTwuB7pysfqbPIOTePux
Zv/tP7JI37l+zgFp/A8JoclXxVvsXSdAGTGgBdwNAb1azoeX2ESpjCYNjHic5mj8
r3INpcR8l13Y8Xb2wPVnmvD82wc0goTPZG5UcVWGmt8+PNEOCMua79eWOGHHGrdC
C6UVFDZW9hGVLVlNfQPU6d34PomzLbhq987IJiRcIpRrDmpGWY7HKZqYGIKA0lit
w6Dvfh1ZB0WzwYKT30W3S/MfdwbM/JRaLN1NUowaBAp+6173tQWcDD/Mj6zVf8N+
pVFaozi8U7pm+VSLv4eXOa4bhuAKda0Tl3I6sf2iDf2cW3KfRPWc8KA1+gftDa7O
XGeWpPhjSy75lfbXruE5vfJVESuQn+LxCO9KAXZ2/ElBkKpL2FGGHghr7KFJ7zd3
dOaLP2iMv6eOmIvG0xbjmxJxwbMI2pDj3iodtO0zm98iLr/WMH7eNFOXAICK5/6G
kMGSFn4cmnI2QD+Qvl8HJoqwP5ko7mHVS88AiJsW9rN886mkofEcebt0nrxDLZiU
FZNJH4l4FTJftdYLptuK6E+/YKRUlptr646/BNdrkNd4fpRIIKOpmjGS9nTVJ2aE
S11svM7dimg7nCjHq+VjVhg9QNyuczYQlyUqek9H0nKRlelTykXMA1sTmrpNd4BP
6fJzAGmz9AUavxAGdY9uC3AkVyllmafIbvvyRYHHRuI345ukGFkmmH8sun1v1Ux0
e3m5ZLioD2Z5ndSXUdkXhTOgmVew7m+0jp/qqUUr1Pi9RbX2J70D7HxGmbdT7eHN
+J/X3sNMf70XEhcSqbSydcwiNDzGzrB4T9MdAVx4IQLO8wsB7l82n4m2dkepDgE5
I+kUEKiMR5en0eit5qWCwzA/JWkW9mUlEHXFGw8tVfpP/QKUT5tFU5orWo/g2i2R
Vr037MdTbb6KerWZbFkiQU3+ABq5yw4A1Y7Dhoxfj/K+1lRhyDRsdDdUPdnnIw6C
DGSiOax4RX+ZrhKOeJML8ELIP7HE9THBWw2IHMjUNmzQHG8pIY5AVj0LgwX6ShJ1
BUNlL8AR/Y773eB6uHCSYxGZ5SPqz4xofKS0R636bAiCadBCHN3qz6KkyygJt2ls
qILfiD/RA75v4+uwUWhzWlj8nwkCUKAM+hKx5J0GDtztJ/LCYHqMY3RZIdCFFZr9
KX7qXcLENiNG70dBYPo8Tau0QAAbtKZX4/gaXPWlo3QhYhSlF7VI1Z9hoX/Lvi/R
U+T3HI22uPeakKpIXNcF8q+gnD446tw5uhI2ejYdKiwV1P/AhLAw+WPCU6hr/8sF
CexnnnrD3N9lffeqXainVttKG7m+KjApSZSla/dsm4OUXN+l4bmeImhVFnTE20xw
JwNA2nud9W1RtEBXk5QOCkm5ngdfZ2Qce4nX+vSMvVZVS2cMcmJddxRIG3zbD27O
JDYZsrBcxfy7OBsCQkySZoMw0CqLJcLUCVPEV+vcyQdkgSMYdzA638CZgeOkWKq9
opz7P56afF70/Y1Wz9cL3dk7CZ6+xas50iT6skA7/D2ueuEBVZ5NZl8TUSJ7OOSh
7EM9RlWQvAA7+4Pi+ymIjg6SEXF8jPhEjIcAqyZFxePFc4esh6s1YX77E7cHj+mW
0k01rFROVviNn9BrDr+5M59q1Bb338NmSRw6vfjbjwoEim2mu0QxVglfuMp+SLkt
d2aV577lF7w8vH0ohFUSgUUp1BpxZ0t98xhGwtw2ZUB4unT4Eos0ZIzADQfO7V7u
URtP0VH6KmWy2mONjLAS/PCPoLNAXpuCvLkbU9Yg1UhP0vZ9TZgasgmdU21fTH1j
tO7fwHkaD4rvmEkzwCormPQB4SBwI/XSfxPJCarb18Oe28guawQv0ZDKex6ywcT0
fFrywtB3SlaOIqe+czI/zYdXarVdunb0BdysPHuM5RQj0JB1g/ggMEDQsiwyHWlH
3WDcjRGP1p7HfcU4Rc+SiSFIJh5mLbw6NIdMwbOHpRjpYd5rIv0uSVHyJjydT+Y1
wezoCFYHaZM1zZ49YlE224hBVK0tCLU+pvIsEPlgmzM+2X/ztkWAZ9dA7tWcERA3
HQne0+8bN/v0fWIDAjZi/jRiH2CSXB2gjBhliGssNSMNMiAfc4y/S+xTueH3KDqO
mqg6TdC/2VDFRfyk3ALPcsXyfnzU7LlDdX7rBTpIh+5rD2MWYM7Qz5VYjhaYHAFI
XWKGmCf8k5wEE64LfbY3/pTnoqOiXQvjrnebnczpkpZENSiUNdlf5Ok5dlF5xVuw
bSuKgkkIvnQgxg6cLcFlauRaB75TOkBaLD9pDPknZQ03PmVre2+tvh8g102s4mOB
1aABOTlcMcWnbUrpYN6xXLbFzKrnLxJYlUYB14rjxRfNkH8cnm09rs92sFu/NR3R
GCuYx71X6iJ3oAsa8okgAChlS28mfEItdGa5hpSHsJRP2T7Oh0WPMStVZYVhecRq
+250gusJfVPujkFJe/OSkcycEJpP/k6uugP60kmXA2lio9dlqB7AIYPpDhftiJDf
c6zjhUHzfj05zjU3uFDV/BSy6Q33nus93xKzBQ/TSNtwiEZdm5DnbsqW90BRbBdD
rj/QBWhpugPrSmibfiAwQRZRViv/SxsjvMiWZOP3k8lNORk8vtmZza1XiLiyZgt2
8y97dLRxkFmyffJrjvPOmNoRkG1jfgAiP7yNC9cItooTxxvjsXAd61kNUnN6xaWv
X03VLGSA+KV5+eX63qEy/IHICZI9JmECRdY2iHOjAIR8ePJEYB6paoEmbFCBDfoT
BYb+/JzlXGKHCRjgNvZ7kUs+WpFmdfw0iZJz54frvrQrV8cXK7TsW8bN/JYQBc3X
z+rElv+1fD8rCoFFcmLMH1+yHhULLa8rsmu8/tn+HD3qGNYhwlF0coJd4zD+OGY4
b7+3B5zG3BRWMeQKZwRm5Zr3yycV5thENDuueZ7jZz2/Ih0mwg0t9LyRrrCh1d1q
YShUo5Sj3AsPjdEd2DrJ/Dhk3ARQwnJNhQD6NLni9+PqSCviuppBQCjnzeJH+ahv
++1Th7KwlOmnI3zM4xdUiVxu6PObi8q/qmgIgiMOm2UA0eObjAsNO1HB6RAw4e8a
i1Z0a8QeX2Zj2v3IIFy1QUIxgnJjXzhbz2d4xmVZsW4XL7jfXEmKu5IyBU9rilwk
/qsNCBtnA6aD1gBsO7M99T5mxzPFPH38iX714XJZdBvfw1F48S4n0rVAnGwZmKJg
38gXtlYPD2jd28xJVZGCl+YmhClfZk3/SoYGkCEt2EPpJ7GK9quLEeL1XU8I/hQ1
BBmVPLS5SONINOSAdSGeTtsNuWcl43QwLFFrUIYU/9P2+buuUt4IRZbnHu8ZI+UX
QQL+A1c4tVdzVs9Fhk2x/G0HZO3bQjt91m9OoWV8ULbLPJjjyYgb7dh7IlIN+LWX
pMTCWzkk5WI8noKGDrAzb6dvgsv9lThzAvgdCQJ6/2/9c4u2VYpExBX8RUAOj6ln
zcaaHsN0ywR6CoCVFmjmSQODKSFXDCqgISQkY+1Lsitm9BqzGHfcCG99wXA9yu4f
NfhR78BuCos2a3d4i88FGrK+QJha5MFZLzfl9SSG/bWbPNEaFUChaPFIt81Q5h+h
k3ZgVguDfyMM2uGgYgoA1JlFEKlfJeQG7Z6+WFhGhT74k8+qDvTGYf4JHdRKnajI
iJM69y+ejFHFBHjH0VSRIEpWCL5hSW4Rv8KdrA8C3Q2ja7fFgyPAFvwIJsdYc+9Q
L5KA9VrjiV3spIXJcNUV8r6lbUTPWMkfKavL3BioOJwYh3fXgw7/3960Tu166SwZ
EKucVZXYINbBNBsUdo5hnP0QxPXRve1lR0jOx0dTgvcdGSuigF19J5xt6OCoEcOF
Kdge5nNsCuug9NnBCVKdiLBKBjDXedERQXwsPMXgg8pZ2eKHq8E7IPw0b8mIXUZN
iS8Sj6hkmxCF/6oGUv1q7Qky9Ifq4Lq5d3yxcDnv0gaBsWWLYOYprWJ+Bvu1J1Sd
mFfBHzsr+HrbSd3bkL26ph/efQcLNSqBLRZXdFiSi57j2Nqh2JGUv5Lzf8l4apdF
0i8rfYsovHC70yb+dRyb9Ud8XCYTGD+89v6W4SG9fd5u9ArR1gNT0wCo109OYXXN
0RM2Dc1b/NryUSYse6y34u2ZeYcrEwOxWXTDDOSRa8i/N+WdXPQGsCKMwvF0/YXM
mstGqMY+RVzVb7QpRhmuskGk0UXvt6jBPDuEhUnvZHDWSWTSenJMA3voPBN2G076
IBbsvMhJeu6f5AnKDWcK4HUzf1TLMcgVf033HPV0r6cvKZr3V9yEWLNd+mCDe+8V
bQsH8AzoAe0+viqn1F6d/xUmugPTLyTVoXao7EC5VOhi57dGCXeTyRiCbagQCxnA
HEuPCzIkpm92+FZeuMxlam06rH9VNJy8jSOlz5UFFXc0VYrWcKCTuWM0JJFAgVcE
U/8d+eKAd65/+zn+BnrekyDEii6GxqUYWzbv0s3LsRSc9AsnW3BPSRa1F3Eqavar
Z9POYzaMx4nHojPNjfCNq6omRJ+gVBJzdwfXEku4PAU+/eP6M6svNtwDZ6kgaKNX
Gy6RQvG1vGy4hv07ZkEBpkGQ6MlyByNwoedKWv5emPk1XJi55eWx3F/dpjRZvZev
ESlgdsoTCYO2olD1LBoXcuMGLNane2VW8nOWddegWXHIVnhrtyfc4mKB43y7pqtV
YZbvCiM45aT58c64HPnQ8l4I9SytR6SWdbtexDP8cRk8v8ga2fnG92CFu27V6Ar4
X9KmmDzogbcqaO/YEcgvlLoQ09K4h/+HSYMZIA+yBsYzVHRjQj8ttChzeGriUTKo
Q3QbdC5Jx3VclOPFDDhXiL4uL2QZ1FBwIlJmIAITWpzQipCC1+j4+4o/Ww+oRDUN
ksCgMSELafLcpuRh0Y9hg20M8j591IfWGMAr/hTBAGxt8B78wz8ty+UlcvxGaYPm
OasBLzrfqPNpLhPCDFKSFkzN66GC3DPhi7qSRjuWipu5SlIFlJxqJ+TZik6VJHoc
n/sdrQDAXmVquv91LYpN6WoFfKsOhjF+NAQSwaLisWwC3ZqhcQwxi0rb+FZviQcL
nrV/THS7FhHTBGw3gNA+7f6NwKVeDKwSQifatbLFRRuBD/pDPC7fMiTRBZ0zZ9Xs
r1UNIUQ3BvJfoXr++RaoyaUIpXfAtVt22ljpedFvB1VUFAVTS/TT3/4jZZ914hPd
5O0tn0Qi5dBbIlAKu/T332Hc9Elbb2qqY0HctKpVDhj84U3VlDuJfKMt+LULhjiq
yiWbliAv+or5zWwyc8lyuCW96b7XgyWTmkSuWjPRwQ1jXB4qdJcy8zFGa7751OI1
rsG8dk8HAXhSRt0rz2vSgFJODXHBg+oVhCl7amc8Uv39y0+0VbjBxdVcdp3uTv05
x09T+O/Www7Bx7jmqrQT/HmAxbHoAe4w9BNrSEHv8RkafswUQTcGmFoZ0JaHgCbO
tvKZ5K/Uz/fDTcGs1buVvkgh5R/AxJE6/jNXGSq4vNApNnH/3rf/TY/ALGyDYJMX
tVkzDH3srFAHmD15DaJ9unvPbXfH/4cLHPDDY68ezIw6BKQ1Cl/t7rPd+7TQ57Z9
FMz6B8T7jZRHFJMgTpgfcfvp+khLqsb23Dz0a/Za0Z2eLVQl8SSx0RX+i2rUn0D+
ZQFZbfIbpMjzDC5lZ8ltJFrL5LxQogK0Q5pMghpiBXUeq0sHRe/iqgpE+e/pr1xk
ALTIU6PFlbCG4W/jBBT8nMg5dh7u7ckSPVr8kCvt1LB38QjKrIYfkKNFQGYFVZ3n
8LQKVRIrKLaEWHNLn8XMqmMlW+EgDyn0ibH2l0WCFwzpuEpeShE5ftYldscBYOLE
uPxaZgL8uDSHhV8v47NQfvuTAdu6tTb/TOwvNtaSgWhzWvuQWxZYd2E8PNjXvqhQ
V98Qs6uyOLviaCmxmNZE+WYIy38MshaDGXGwlV1bDdOp8+BRphF/VBnSQSVviv1s
qJxouXxCUlWmrUkwSmYyXGr1ngKxkYyA6Tl1Bq0BsENDUDCqLqrogda3Zz/n/PhZ
OUEV1JEf+b7YA7aYaMjIxcaTvfQvyHEA6iWs8NMm0ru8yFGaOVMyJsJ8vR0BuDeI
q5h36Yx4KwkIWXQ3EFRzPSmFRCfaokXKfgdtka/HLy3pXj+r2+pzh8XbM/MHZ48R
GA/pSYyHn8JocbnmhvWQGx7HqqAfr54fQqQCETI3FMNnDM88KsoVOOwCPmXPfJ9E
MEC1FbWmGdtro/yXPgerNyFTsyjkpWTJJW//tUhKV11pW8lF+TQpJRIqI8ot8sdh
rdBJxNagJTqNHY1kEQHvdM3jzntx6sEcMOkLle8sozquP8b9C1R5earKgUM7vZPk
fVyxq1Dd7pk7Gu9SanYcExJmximCqi6PDmVwoBpN0xwKmf9UkP0Fc618Tfzze+OA
8io6bWgHHR6E5UEVAY/5LXDcAWSXxhE3/oRsCpVBbweBkFRPAmm1Iv2PBorEVxS6
ClJQ6w7Q3GpwkVDlJ4uMjDx9u4UWF1O2MKhV3xAKH3bzXsl61EGGmrYVpZbpeqHS
77daAfeWMV2rtpTax8x5W9gkq0whzmvPx+6KwG1a1EQmXPpb7Rpr5S7fxVt1pj+d
1R3dtcl1wYMq0w2+pMst3xQifVyaJSmyjPvnK/rVaLR/vi/vHe17VM0aaduTGD+T
CJdsuS4cABiJnezMqW+Ec/jfdzjZMgNf8b/oGMmqqS5YP3Und0zLIV2hplEa3ifR
DgWYssiD+T1P3cil+78PEQQkL6vMPCzrkaz9o2moY0Px/o8U0lQ96rEujBeWWcwL
RXRzxMmgicmRKSfF6OPP6WGS+vcBg6KMi6CYK1Sb9sShKl4uqiqWhKJ9D9nEN/Bc
/hMCPZKF/gAF/C0DV0nLrtBAVcM4XdBeNKMF/zIlXQt+S2j3wSnAdCUc1mBM0NdU
VbIGPDULHTigIovNIxk+4dSeiI7o6MvPan2+cfckAOvyxOuzyYqPsf6k3STwXNyi
EvwEV6I2+2581wzQS0O5MxmjyZJGJo1/+BNBTFjNUHpsok/9TrJYSdJkcDiFO7iN
0iXp2kwwdwL8tclxZMZwUBlq5ACEXt4OS90NFp3h7DIRJ2B5JMwlueLoI0+LDQP0
vWstakUug0KWBjY2Eztu6uJUn2vuA/NdoSK06YwBC5jhCJXY9pWM1e7NUJ8OTnIh
ANdIsSTN/gTlqlX3wRnGbZgbwaSkXu1gCNDlo+iO12pCiz569mkngHX+0ErOZ1nd
MIzT5Zkf/hj7Vct2hwTuG7Wrut/jRB7eAHcRAOMLCpvt4oAJxZSFgumpHhKxooAi
4TsYdI7TWx1p2S6GhpplSvoKmibZvMDUJI9LLw2kN3hWqynP0u417c02YsiwZJaJ
a+nFTyxxpRJr8wGs55CnMN1q2vjZgaZeO4Q7NbnG03zj5JiJLGYHM/TZPiyajRQJ
kLHdrU2XQDz0GclbEXpjoSrdp68SytP7RxdmBIz9+c+3RQtKbVpAaeWmr6Tam7n+
pP29KEbsek8muLzQkeQX6cfZ8PdNs/4ABRt24H3z6UXX37lO6JHNHBxtvJi2Nv9q
sVkNwf4gp8UFUMpNBu9Xi9a85UUroXVt00cClUXgTexzY0FDk15aUSo91Pb/LM7Z
JQh09MJLuRSR9OLyRwjDDn319mMtypdxxzF9Ain3+dqzYSwqcoc/539gAQrLmUCH
J9PG+BlTJmvNf17JQnyKUL6slIV7Fck9t2j/te4YKS9he7SxaX3j5L4XXAZZ8nUQ
y1OpcqtnewtgL6e/5jJAeSPOT8mY8syIXYVfNWtv/u50YcD2nPTR1OWnoAZOXnVT
tn6bt5nwBAFZr61Yel9DgxPKqTu/NZqqfXFfFGlYDkIXeydIVbxmXdnKYixCDL47
xdGH0LduE+Lipb5v/R37sVjZ1bqJHl4jyhQlsYZDIIOA/PrGz5ENPXzoWwJVW4lN
7m0Mmvn6G+PvuEe9By0CUG6vay3lYlC5zS4p1z9HTebohCW8pWYBqbpsDhdssKN6
bWYL1x3v+QqHwyLyUarli1tY2txiCyK23oI0wYnEPcMzjN7199ao09N1NE56OLja
HYEicf/5/aa/3WGmvFmnfZP4ixBzMHkpWbLyzNzoCEhUSafqZGdOouhzCYYRnrNw
o3Kkya0MWQMVVOz23Qb/LH3HksRtnTtQ6PPGAOtz4gpYSibmeFUg7V61ePgmhQj9
LZPYQyDaOyCbr9qrhpGaR3GglHabDVPgJxQKQKuF4eTK5lMCftBFZnoqICmTnufW
fXdWybz5nVUl3DswxT1RttXAZDaMZW1hWMF1miCMQehfbf9tHkGTQBveLsttOKka
blGGM0U5VPigKeHeglK0wr3TvnvRrkviNhCzG321S28v0mKZbBJ70zU6KzUj0+0i
i9eu1JHkJ+waVowJ4xvoQs3IojunoagIBZJGenKBKascuBeiG6qL6RvnDc34XrmG
fOXdPNB6U8d+GtEGGxnocTlc/npF4D1b6kWMOwQzj2OrnYrGHEhYs6W2VUqCMjST
VIlLA8lP08HMBqXnxKbzwi2peVPhU02g5K3xKFfEuG/VgtCBaiw/1q0MuLAnJz9M
Mr3IA1W+jIk6y1CCJMCPqAnP3Ahi3Snw+oGuaXZnUxwnLc4TFAwQcOL0ABQ0TLz4
9qrT9WJnp54Rk3qoYMHTM4tuBOBnQjle4MGP5EgOGhfp5u++IjALqNfZkemlPq6R
dRiFIc4Wa3NXGBAW8YlX8hZ+wb6/QjRk/CXQpMoWmZvbGRnBPnr50vPhZcOLcCy6
fuKuuuwyETz60UtWcosQ8aRwR2p8rkrQkg489T2N3zh8pcSUxaIlQ/tRZVH1cb9v
jme47XVaK2wrxxIJ1M1hUUHXcgq/VcrhXuyp7pPBaMf5CJLpE/b6SD9TQm7SjknX
hwzuAxs8Gvej+a2232YVD2aWq8rNa2o3OG2ojAwQDYO92HseWvC3X4uvWjuURYgv
+t1kzXmdy5QOFonnafwAivgWX0sq/JAFG79llV610xmsUw9IdBE7lZkYtNSAiX2v
KeSoYHzlax9voFMTokSFecTD3pKerPUWrt4HYf9BUUw16IWrzeBwDZqdziIXnt75
CF9qsu555Hf2QfUkzLsy4PjGpYm+FNSLI+51CLpX26pY/3sXPjQgUC9lxyJ6/4q7
L6m/ZieRVfpzBX1HEH5t/NqdJHHWzM+wnPPErz9YnLLoxmpWmqBysoH9K+fEtsEA
pFxh9rIfKsm3OrsaNhkk5rIgult2ER+Jrs+fwKHIiyRXgVY7Ldx5yNbveg1h29ya
vST21AwzFYtMGhxyW79GnaKMHwFuDqZWZmMNrWeb/zFaid0EtefszeGdkp9TfZ77
MwbxAjSJevK9KfjEqwP2gG6W7e6saSwKyObWNl4+T4XZ8e+1Ft50D8xCHd8m/YB7
UETItulUdqULOQI0dHo+ZfiFvEh9G7mqOhZlXZ4eBuL+F7rc26ZZpGHYa/oO6Vkc
Rl1ZIsE8VslnToDDFeL88faHhwn/YdZZnJPrU73OBNmssfbsrhOJp3K1Mgr1BQRQ
HEHuo5QiwSQipelHe+Gi9i8p2LGPtHG/yTtla62LxwlgPO2H82FFFrhBW9eJspfh
4jN+au7qHsedFQU6ib7HTXc6g/X3qm11+x7ylQvMr4w/Aws0B6q2MMDuMNeZ27M8
W+r1wOMrS7ZLov8EL4p/kwSD3KYGsqn99D7efb8r+qOj+8srY3kp8h/Fr/Sw8YBc
+3PxAPz1Uh77Fp92yt88oDuiv4fyjEd5fjDP9p8STZcnq49XKcnGA23Z9SBP5YCB
AWNZPynC3mNPz1rk0XNk44KQZhnEvjnJhC8pI6odq76T2U92UG5xJJDmA1Cc/Iiq
x29kzWZTEfmoWfoo5nanquDP+XMXBC/MlzrGJigAAhliP3l/TvnFgeoJSIeeZaDz
ReQ9zcSq9WbGui+5usqmF1EwO9xjVyfryRiNoyX0io35UDtUYSj4x06fHUrSQjPh
cKF5ntUmRyg8UUPxHZ8MSu9zL0wvElwDnnyi7/56BgdZYkzir6FmkR1ApFOQ94eI
pKmDbnVq7R6Z6E2WJKbc9MZHiaJQZ7aVNbzYX6lBms4PObKshHfbB7bjpdP9XiPZ
PZ+iD2DhShfxdcZf/3J1Gp3MacdnNc5sJh2IaUPQOklXuXPcWdFUQMhCBcFzFYUR
Edjs1Jl5fLhs7rgwWk2b28az4liKD6MQtoq39KYNednWM4T+ytEr+OsAOqg38+Sn
40MHTaE/aIN4ipWVVsnKr65PADLm3mmUKlntzWYieQ1zp//VOQaaePGZGlQ+Q/f/
jNYZYjbyuiluKgsFp4nqDwILKccLi7A82EPxtyJyOd3wJ8yxhMmM+r+hcXUHUEVN
Hd8ccUHyw43PovlHPzvxqkMlv3Houem3u3w5NVnfB3L+B7Nwh8qvH+m+EtV/KjPU
WlmVEgsTAWjlAjqjlX2OAmnKcAC8+JZW2ZcSplEaZ00yCT4raS0SDZBI+PbSs/jP
mp/uUxa91rU44juj9/ZmE+sMyjK8kA8/bL4o1BZxcoRp0y8bjVD3fgcChUTdNodS
41L6Swa/xthtOnF0BFOTT8oB9fM3cbjF+0sRrfzqLpVJefreS2UNLsEQt5+yo/XW
L0fgI/yk/qdYviNq808HjHsqqnWMU3x5I63gucx9WoQsRz5Bhr0a8loCvwT5hma/
ysWPtWzK/7Cu0p4YIUR1VFZ2QFMAVCGtSi8ufDwkOJZDnbnU6H4Bec29eNrjDq3r
kC8j9XRpvWx2/EctkDpQneYzE5Cv/m2h1dLDaMDOpHWMH5lpdta0OzjQznWC1Q6A
L9A6ALZ4flbCh7tMR4ODUKUi3f2SS75kcUXZoaM89elTB9PnvGQJWvZsslyv1dw8
hVmfTLvNneeeoqdfxtYRWaCzm2bGaDN8fXBR4GBOkH/o/xG9HvyH0NCjy7SR+AjP
wck3SwZJ9VdrsIUXAFBlE3A6jGSV+ea74CRltEfTRcOsWohbi64QcMsDO5bqisSO
5rXZRyamU74xaikBi9OF3gbuv1F1/4qxYBNcqkZgZ+q7w0gzf9fiKmcGc4982DKp
2airMHAft2RvHCUDj9YvNzcmdCtA+JBALzfoiZPFnxr0E7vHN2XB+8swZiEoAaPP
NCDmiO8r90TlcViciFK/MdiV8ibpmiOPBkC67NinvmyU1hU+1CchjP6OnF5Tu8Nc
uV1gjNtllIbNykZxnOP0BW8mpwaaHNTMU9JgM8u5jsaRpOhwEmNXzCi4X93UHKOt
yYeAeS3YLWYCdfj/x3faSCC6lfkBT6oGi1eOZtLbF3kWbXOHD3aEGLYAjNQ7gnTH
hHqB/kOS8HHpX/FoAKMGFEL5V1/xfnqndLv563Hw3K8jAMjCrCxSElA+F50vagqL
knM6RT6snfRApBCCtuyYCgySe+vSadItd79USf18pe36/jHdN0gvY+BhP+Rn1NYr
Kj34OD6q8oNP0cYKHJApvEbXkJ8LpegVUFyiX7nkTVh6XR7l07flo4Cv+PfCNjPP
E+z2ycuSprCxS/AxkqfK9Syj8uto84aPMBRrZqvrE4LQChh3Rndnx+MocXnIAaH6
AyRy/GqEuzvbQJGhHlNhud5gEE22dgFhlVqswN1AlKWMAO2jA+cpY+iku6dXME9F
Jiw+kMYPm0WwySqRWtW+ZiXpIdDzMZedURidzrEcS1yY/KZOoxllI9vzhINlu9K1
ewDV7/CQosu1giAIWcNJyv7ZcGqEanSFKZd3WoAXHgT/BKxwigjkszaMzb2PM0Xw
gS0rSStBg3ocy0+a7Cg59g4cvmpSh6gPfi6Mk42z8/KmAe3I77bCXv/dDmY7LSlm
2kKt0sDfV7w8eBiuIIrUh+NuNI3Emvp3jlypZeYFvcwK+dEa5B3J/DZVpU3/DpHj
5K9QOmV3NWEA3cFz6z8ZM1ms8WThhJeGmfGmHQkclf8sq5LPk2tFcEmzlZZ3zjXI
XMXfV2J1jQ3/TSlEqUznLJCFkJcFwW/QC4pixMmzm+eJQ1NuyOh67n+N+p7RT0WH
iJRd0xN2bDu1ZiQYthNmL2i5UFj170Joyn9hV8rhet1GmIXTJAE9DvDNkrqCHGQB
fOlNew5BfFQelp9HwBeD2+gYw4yA03Oyqq7bV0DltK+O4txiEfcKprNblcsX98KT
CpTRCF+NZEYX4wmMVRocvuNl0M1NFC4+StikNt40Kg+yGQq7LvLOFo+YySfjr88w
yOTQr9xgfZViUz02R6KVYc19KMSsD1GLujLcwYyJwQWLhI8WdUoKzQuQCB21q+ug
mpBYMpPaTIWa2UfM1r5M11X5DxwHeQFNAQtk6Bja7J941JhdN7qaENPNqKkGGXyF
W9ntT7VD85pYtqWMjgNontPvdRcXYzs0NT45wT4+x8CFbRnip7ATpwtBBRYUE4tk
6wfr0Ebka+qLkWd3xbkzD2aVCwMzfiwItNlhR+zVgNBHMyXVMdL45H3bW8NfySrJ
CrpZ2IljBdOk5l37KltsPhiePCVX5mr4DfwqQ+b80R2pDZoPgNk9WHwCPFFwjVjH
aJRpzS8+AfCM4hpPfNCsXsirL13+eIjhgtk1NJ8vEHp2KGVmS1p1I/fw0thB7see
Lk3hF39HgAePPCEV10jwuA85bEXXndcso3HSoncGpvBk5//O1rZzw73ZKzqZpqpC
WI4D1wmm4AjQyqyNsefM7SPBlx3nw/Nhz1rpP0uhwbiQeSKOh6ghHzCOc9dqfXzg
/cxQGhqQ6y09xpqwM9q1aL2Pvt5XoOV+6tFeytWdnGgNZCV+nAekwDvHfjscHyi3
TE+ifo6dwSfnU+FoU2cr6xqOiwsl45wAxPmckRBAHNkeFyfA/EudTehau4wWeWsj
edVzd3xM4nsNe/+5j9bpCwDfbda1s+b5le9cg0Az/Y9B+okeTg/023OakNvZ3bHl
TIb7dc7zHXovu3Te+CzG+Je1vf9oaSlga9P60W8pq5AyRUZoJOQ+LWWIUnWYuSAU
WvRDiWY3343St6U5ckk1zoEPwgHSCssw8n3U/H/ucah/91yXdVIeV7GgMBZ5n31y
cnV5zSxNZxTCdMpe9lKEEhyL2a4Ng22AvR1NNydzqvg20/mMi/Ff84jnAf3dGwtL
EoT/KQWm01K3STPtPf4/6yxzDhvPHLMV4d8288HF7VxAZ1wzaoP7bQRHO6EFTF3J
WE5B3wnD1QIa4/y8eW2A9GJS+SRsyHm/osSQ8Sy8cFyC21bGEVTHSc9hauacaDS2
xbKqyToixJFgV9A+hkv6BK12ywZwPBGOv8DX2jaByhpp5e47SprRVDj4yT79bVHY
63Uko4CgdlzbvLmVoE86Y5eObW/nVf0Lg/agPzQ5wsagJBzPVpQRV64ScNFyOgJk
fAXZTtQlWsPeGh1T5H5Nu2N+pSUCb6ERBLhIc2JvTYA8+YT//p5iWHQzy6bcmKfk
v1HymRy1ElFJIxc3PR1JPY0A3+T74aXV3PPE793MKw0J4vDMdrGxR0YmXOCne/Hw
PFp5b10wwxaGGdM+hEPWkLT4H2njtTsKa4Z3CNAIEvwp2suOUqniH6f60izd8zx3
f5Unjia/dYvdLb6EhEShekgjnpWi0mVA+jW+L85BZ7j9g4uul7hXbbe2P85nJiK9
J0+EYCuPvLKHXuQCb4hmVk9w2dQyuUAy7hTIse4jUI4AYaXN8Al1RRzEc730TUwe
T3/pfIrtshNRFPFbb/Hv+YhQ9hDoJFMQPlc3wda4ILTyisRk5B18Taoib1r5kv9/
05mlkXVDf7o5RzdhMyhlFYn2nAWTZ26jL88pQ9Tyx1oXKrJjVi9/kC18kHqRDorH
4hblEiD/VlDiic735cDFmWrG1KKrz8T5maMHKE8P09N/janiXeU4vZFa6t4yJmWu
4h+Q9hFu3kbDB+PHpggAgHyAtGzLvo/hV0orCFaH6y2k1wtqwuSFST/yz8TKFnem
1otCtTt0dJpsev2CvYBwEMizklW/aM1Z6rR8mPAV/Nq8kWN526y5h0qdnv2kemV0
i2Gr6XEK4tkgibsLS+MqlULwaAyFE+O82uw8sirHz4/yLx0RMARJgFIYeYc69k+u
voOTriErpoFS4Wbed1tyjfA6lweEAT7H9viyVl9coQBJ6JWqW4vi5dCCrto1L8cE
ZYivc16Em5hw8Ra7Ek0+tdkwuFHI4AysYHq6gqC82VwiB41M8pE7p6RJ+mRfk174
vLaJqXEvsWL2KYkTCdoTpMLfRztF3Hy7YWKQw7y2eGd7qRmdE7VgFI0b1GPjqzEi
5rDbGaFspmXLjfF8LyqXjNWEOJYaQht//78Jltt8CfLrjtRHWx7n1ks/gPFhP9vl
g5TCk/mJaweylG0qaZNFR6DnoYqKmL2HPd/h300wzmi7aFmAqJ+TEa97pkMfiT5+
yPdGv0W9OxVjaXZRNoUKb6WpOkdkIdM7hmfNbNwNolT6E7+nY8oxF0BqhvZ9EwyS
1d52BAYVBw7GBA8EUKdPkO+Asmp6tq05+zi62fA1HEMd+pSdUJzgRC4WO/QjksTO
zyleetb/N/KFclzCwx8AdGefczBq4SULS34sjMQZ/TGhISef2Hmq4VrWeEzGVpnq
6tPp0nZuleRW4OuPbA7gUYPguCAv6Y+r0qOZp3T6ApjPxrQzo/iYOCzYOms6I8yh
EmOZ800wZKAJm2wiZYvgMqm3LjZA42kHShDMpf561uAAvhxYg++N0O3LvCCiBXpE
CLceoKcDxokUkOfJOT27VJJwPeNpZCPsBZov8K5M69+wv5jRNjZIbTWtx6YGKKre
6JGzBBIYfZK4/grfV27Hy4VyBcL/Yh4ZjsbJKD336dildti/qRbWhG43fgSpwsS2
mdh2TeOTkKVDZKKMz5220Dl4f1oTZN31gczklcu2T8cqHjKQiYD7bEsTd/Gcg8z1
3PiZcw244iD2/ZxLps6g1oBSRBJ8AbMt7/9MWrk8rOFHaZsbkwZMV849RULFIx2I
mGl8BXBGf6ZDQxAqfMIiJD8z7+RtbiCe/uGtDDSSTn++bnLLucWgtHVIkZI7IpZB
6aPKsMO/qO7Z1gNraHbXnESlYnzFfbh319oDMvac7LjGRI6OEE/juM4eqYJb+aOp
5R4u538CuXm3Mcu/yDrPk/lGPOOdjjaXDDPSWYAg43wZOuelXtA0vj4j00cpbtD/
vPhDmrhnerhlBjTRH2IpK4+UnQzD4Oj3eXwiqwcK6OqyB/PW3xdWYN5tPzuVzT21
ijsNjNjyj465K/wfPUssdmEYJalz8ogy2pMv1UDiQyYo5zZY6cIUPoontaugHLM8
/0mK6fZCH/suuMYO0RUObJk95ZE6Bjl0ThfHjrXyOxZObfJzN67WJMJXIPBNzlru
vsc98EQJnMQstj7zfC+Jv7EBeWMfqg1A+o4lz6PhVvHAlA1Ru3wG+mgn4FqjeNnO
BtRdOJBXU92T+HzG/NZC/77EknSbWg5EzNlxLf4r0wWco5tLHBYPPBEinFqFIRAw
g5CuB7qttaMPCDr1EGej8lvGA5WKh6qsEC0uPAe351VZR9ZAXsppAQqxLEd3Vb82
R//B3CjFag65aVkV+VP/UiNc+wYl5cn5iS6bdFC7PZIiaHhkHbsj5kIazZmktob3
iskBZVMdwXX2XfO5JZ8gdtu2DBpmvJjTYhjgd0C7vxfyYIbXFxoSE92KCDLwhsB1
2F9wGY38zJ1tszOV6D9LYx8D58i4k48HKNYqhBscWnSjcLHzEhkOvJ7I62SqKk6x
T2MZ8+FwSmzM15cE8pojYkf5djmNI/DkbP3OJOVqHUpLs+YwUrkm+kG+nmNSltuH
08Ge+qzWBRGqygsrd4QZaYX/gQwijIti/+6jv2yoGlsNPE5+I7UMwZ2ltCOsKwhl
i7nOjNAeNP9/DKWyKda3lHHmaGd8mAzI41kfdHeW3rTaCvTofk5B6a2in95li+zo
A60a9OpW60RjfD6R8yfOkBcX2ye4TbIi3fe4P6+DRrih+tFhyZqlzwRbmJHDyZBl
r5dgjS1ShdAQybl4xQQSeWVtj5YW1qjM/kcvvFzm6+rkS74vTj3hd1IEPmqByYz1
LBayXioNSdV2/BkR4QtIELypxoN/i3o4FWup0RMGDj6kAgpyXsPEjN+0GDiNdPvL
D86Yvnq5dHUu11Mf7ZzqLVfMSDzu8+P/Fd/F59CnsmK/m2atFjq/nh/5cl8Yw8Nx
SdMqgB4P4WaKWLIQ6Ym866I4dValYk/dF6X09LMZ7+2y5FlkuoQNwp/d4v8u8oHj
hz1yAlFF/NnZCGeELxdTFd9u4/GSojE/6YHfmhTncC1oGo+JK3+MAYSVreKhWlRB
UcDtZNO078zMzPTGKby3Xo0+7L8Wt3GMMWnfSCFk7hfRuj3e0IhPS1t3G2jDl9M7
XflkBSnJipoGI01wph07c4b5flqO6+Nt1IspumpZY6d7SkGsmTm05a4lHgO+jDEc
kt+KTLyJzNTmNo7JSYjzQX949uDJK1tXhH7AcCloJmWCAx1wYyskk2kUb7pgj0HX
D/5g/4qK4oD4sCh6oYKuL7rndhN4r4TA2M2+dgKF0SN/Fct6BLXTqX82GjHz2+Te
/weg1T3K30OS1sUwXzVx8eEwDy1t0CKicnnKaQeNUxEEmRzGmMleBNrpkb7fBezf
+gqujG1FrAtpwMw/8hjnkWPX2r9rQr484JjRPsik/z8iIoXBx4oPmzlOXdukMqds
KexB7DAJEIVUdmnxYoRzAhhS1kr9v0NdAS5r2wVIC0QxfaAX1J8qZ/ofaC/99KT9
TxnUVHiy5/b6w6aq9OREEUMm0snycZ0lu4EyqiWslOoCPAtHou3I4jooanoLUA05
/p8Ndceqv/VOoHArUT9XRzJbecxC81S6xmZwTtgVQzbMe/2Wdvoq1LRETpoqaaPn
5/TOvuOQrhgXjSBXDMwr962QlJXKGQuqnA8b5NLKio+1YtKVPAKzjLW46aByDqei
oxxnGJcLysYpxoGwNU7N9CDK+PMU15a3SO/jaIZzHm7aXcthRZ/DA6ongUmqJCGa
xnGAHuWGSg5VCjkpv1T3UsXZHbVw59sdjKaXmq6J1QINkTFk1SgX5C4iGE1lyyWT
mpJ2PdiZZhm2Bp07+PwLuD3IbLUoY4UNlQduDMDpyeLKZuiuwEbejd7A2ehuxkvD
wYJfMW9TPqIE7ORksrd24yYN6Zo3HI7w/gFAc2YjDMf9kq7oVPHbrMMMU7IcrTlk
grkD3PSVymHjuQD0V4La50oNPw3HrEyda0KNCUtrpJxDS5JFBzMFYEKyZlxaTCiA
b+tQIZAdYL6fvGIx3lnsxE8DcfP0mm1VrbSRnQLrSJR7m3hr9eqs7RBAJ802lo+i
KPjtUdQe+ifhGsJ0BuoCg8aCCpiWDqjLmErnFZNPDCcqSvJMlGNi5IQOQokxvE+X
jTE4HxW43OkIfgO9o/vHR7g6LsSVWobLezhEwKFVvAdPc4lNdK+xX+LzyJAYZzEU
dTPYxhvc0D65a8L7cuWdgGkt3Dvp3pX4FZooCfEZ4OAjUEei8Z7ZsJYU4bLkeU6B
fetAaLYAAh7iLG6+N9f2vyMCkWcUnn9jjIodYHJDu43NEV4ZurVHCrX+oi/VKwJQ
`protect end_protected