`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
dYVY1GBMsK1ODCn3ZUp8SoAWP8Fvt20jOclKciHf7Ysn2OlvHpNHbXI7BFbSBeZ8
c0HSNxtSIQSCmTTcVbiOe5bNYdnShY74EmVDlUagwaODhK9Urx30VHPfg7K0Q8Dj
u4EuL8LzGtWyNpPuuYUPfH/EWWJz8j2B3GlAugKl7fR1RciktYEXyNArDzj2i2Lo
icoQhkynNgC7v9DkMLR1BxAwtrFrckccZalCrbzlnjwD/DOLPtfjLaczesJPkKoa
xZJUnnMJHmZHdGCWDxS1eicDF7kXXzsE1BA2jAX7HQtg/mw+vmEQXKqvkKy9tRtW
yhUEHOXSIVFkC6gJ+buK9Q==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="SgR4h9hEc61j3UcDg7JP89NUc7gPf41F4aolx7zbZ/Y="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
PcTZf+e633x3tw5Pd+98Hvg8K8pEx1TP/UFyHup9OvIvZyp7VdJ/eQ7Czw0TCb/d
NGL0fQmqipTyP1VBR/CwCDPv8pUq9mWdoIhPzGBVMq1ZfAiLygNMWUwFu0/xPfyw
rAKvJfKF1tLDCsja4oREz1+w00FDmJ2gsQcbY/9d4Lw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="fB5pBzxyhRsqq3gFtq6qZ5Drx26WwP+GzJuJsgJq2oo="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 200784 )
`protect data_block
Pw0LuTSwA3gmWF21w7rVYBcj97hqvAcf4dxm1w8M8xOO9V5Zp53fD6281Uk66by2
V+2le3pjRQ4JkfVvu0vvltrqFdWvBln4SM9xPIyOvOgxR9dZ/mACNvSM4sNQA0B/
fX7fi3PTNZC9xbat5PE3y62ZNSnndh/KjPp3L8rurN2Fvb5/ju8YunzH8nBf9dL8
xfKf4bgt9Rn7oDR4OmbwoLPF8RuH3e/ScnY0TVcS98+dF2mPhPBQdjcO5DPO24MP
DRRvnyvqXbJ8j3b5QwH0O39ToHKS+ObUeDlLRdf1Hm6zK9JU3h3BSI4m4NlXFuSj
XntW/OOcfYjMCJmnRNex7/Tf6l1+DC6YRTkbCn7ymCFKQA26g8peS6wh6k7zJDq+
uWNhRRv9bW9b6aFrBXXoJtplXceM2WVfOAgVVJT8UStD3GbRsiiaB+/3w44mnkRX
LHPHfqua/lYC6qkCwSjKoF2dt+o5Xq8pTiFIBmYIXvDF5hbX5ACjAv6enwMY69tn
kq6FYjprgdjQeTzZCM5NJaISMoyJiMkOYdPZWBITzIdN0meXMuPv2wNc1Kd9r9bs
710hh4TOEE1/BOec7wv1+iEyWzA9QhCXQVTFBMI4EE0yLGJ4JbETGDxnceXQczTC
0dDvU6MPCkBKBWwIZfdCAhBFqoITcmAhxf+TCjvN+/2eKJd6eUiFaeRjjxx2SApn
gJywFiypOhxX8jU7P95LQ5esBraCNGAekYPwhhPSKJHsJ2l5o3uyc9QKmcdQJxP2
foYMa7nLmCyfA8nr0Q9rSyPnDAzrxFxdWScUoeY5brF1l9xvw2FGYKVHrIk9APYD
FvjT8cXKZa0FrflaxMdopdE+s6mpZby7BWPXJbm60OtcyR9qx2qbScgBA2O40X/s
R3A3YLeRtWOWbbMevFIkpzrmDWMOP0NogBT0tRJktVFoV2h9h6jak5ABiDjkjrFu
0pA9BafJS8DDFcnobuuNPbo+eq3Q2JvRpZZedd/Vq7DqG+Hl7Wm5gsSjWm4yDpxD
DaLLPYRxbYlqk+5w0OIP84fuR93yIEJSpUr3D8hCUkEx9hyB4F01LDiT1Dl5CM6N
BNbaM9vVWPBt55TH9NqpeykhgyWpLZK7qKCeOg8zODp6BRyGo64t0UnA0q/Nvv0l
D3R353wvq4LT9mA2jCjFyAaPmHJN9Sb249JstIuh0ci4sACUPv7tBKqteiWx8s2+
XV3Je2tFhJMI+wCKiq+ZjpXF3IkQwNbHQ4b1RIsNRv+wKkLA8TIUsWtjRNOdIDNp
PiybBQK2R6mEHueseVrTJGtOWPmwima7LT7l+pJXrLmVhSL4oRpNbOjW/rLX8Pd4
61ugBPW7Pwujzii7h/k3AgymSFhhlLCZAeRU8vpxgNnV6U42Fti5nN/PeNRv3xHo
9A9r8GqVHHsHEb+dmX4FlVG4uEGeebKjy18ceHFQEjtzwrOQRDpZ/iq7aAw5uHoJ
NeRSwke7WgNgmBYWiJob6zPymxf/cK3grnb1/fLx19fx9AngggVpQlUx0btHidgE
tVXewWky6XLSz7N5E50GKPBMpiXtSPmpvUsa2vIXsNZTOwKT1lZwwCiSyQl6pj1B
OcYMwtzGp0YXYXGaKvyJlSIxAMMTQzkaycBjgdEbWN+xm7gtDfCo/xRl1rmWbZxs
V5Ix7Fg6f5dGAFK6gA5gYagCHUpgE4FEYRdFX1I8/vk40x0EYc3yb+trwme1TKna
ZauKQe9/+44UCoktWFNqUCW8/13LxG8NSS4dsvM9PfmoLXVVPDsQd1toPyFgDNxd
AjdJpdrJnrUifFwYL+SxgpoowQjSH4La0ynHMsrPIUG5YnizfodUcNj33BggQ3F3
g3nFnXWdmJ9AcKG/Zt07ShtqVDmS3+iLWnzqLVSpXq8/qixRFf24kSfP77SNvn2J
awRJBhnvtjJFTwAWjU1CfwGe4g7OEnAd7o4MYjiGhsyETULE8RLuSkEx/PIcFMKM
v8sAJQawG9NUIU53EIaKjQ4M/P/czi3j/5uW/s5JmZXLmTuyfPkhp2O3UQuYnizU
ZdViz99agBrXM2kJDePBM8r6IDLDN8VxMqfjFbvVJ32Ce090cVmlo0UomVxV5LTX
d7JcVOQJzZdB9/nbiBYelLGAtBD13BYhnOSrT0RkmxCQFZ0QbpSor+Tox/JB2qgc
1IU8h0w5T0E47UqWFpAFjBrFrgDBy+nz+LRBr1FuKq7I5ly7NLI/WR4Sslfn4p10
wyBlPgtyRlaCCKwd3O7N1znBRd48lUTTmdL9HkF5I9gwTxiAhHDIOjfH+ByZr90b
8efv4PXOczFRciOTIEhnOFxduH3i4kEqK3O3t9i1sOLfqA3u5R5oy+KpDP5RT0+e
IJQq4BsJvKgEpIW+tIXxJnZ6etj4Oet1r6hZSg/+7QVdajZ5spaKt9wo5kkTM7i1
l8VuOOI39gkcq9PQPpo8gzptGqok0eVUaYVQtvf+iH2pps/lR4+OM+5qux9w+Bw1
fQvZCpNR2xUW4Q7mAhZGT7dN1VgcDPPwK1PDarU16c3AeuWoaq/jFtXJtGXa0LI+
+fTsdKbUXaZpY8tab2n9kEYSPEgzf5GDyhF5uvwpqU3QrmxKxXKVTst2ZeRq2f22
3DXCSvlJhO3haA+Vy8SU5QYK+01E1gM5tKtGlztONqjiVgb604SBUHNgpMVqBk5d
6x2VwJEfth3YWZB1VPO5Eoyu+ndigEtPbaDxtM7EP5+ZfRLc4IepXrD90SNaBLiW
1+CbWyuut4RjFGs6mDkuzf4zFe1clr9hmK1X034pDf7tYvCIEwz9ZGY0QlnBCloX
Jm5PZ49ILyNuv0yJunaeis7870bO0gPjF1SSa4ax9kYGm9aOxL71F91P76ic70JQ
6w4LOLmQ7wD0s09EiW8Tsc+XVa/Y4UMECxYUTFwmW1O73a/wmkF5oofDtkl1vv8a
toPevIwkcVQPiuFNlIYJvqbsVvCCcp+2c0j84A03gXnTnF68Q4y43NfHF6OwpCcf
N+3z/NrFA2bHO4Qn/dzQKQzFfpe+meUmlIlzBME1CpRlZ09eTuYz59xg2NNIxknP
Gyul95tr47D/eGUGK8H5o85mYyUOMRVUVeGLYz9ECH6lUELg/32lZ+BoF0mYqta5
hHVvXhL0vOr11DsUdmPnI+UgArNLR/6DI93hC/BlvkLWv+GmPGWroPfV2vNrg+/Y
vYHUQZehHbN2PgptOjMRWHMJn9Moik9SZIUfI2bwJhUVM4GRfwyv9u2Tldwln7pK
hNvUZp96/uqJHL4mAKriIleUCCYJ/shbPyXxOODrlV93EIv7gLw2cvCG/SlcRh4H
p8w1W/aqFXJOG6/R2CtZf16omw3wyzH1ytB1mDremKA83tLA8YfFQ7aoh58yjajj
Zi+7yS7cweaEHgghdJOn27nMHY3PTPrPcH9BREkdzWiUcZxwB/IeYQkaYgH4O8JU
Mv1cooLCQJM61phZpj6zE8p+URi4N/RktlRLibJ5Jnaxc1zkS4VAfUWdUjGim6SL
cADEN8Qx6pHZ5odBDEtRf0nC0K/7vBJoOJT5zTi1PEpoDINrKq7pDUmqKYRp+/Ws
h5KWvaccb80cfNVwzIO6GkpxB+Bymu1muZJZwNBXoP33HfrbFz98jFYfyfiFoixl
UX18rGNHAf3cHLOHeQcCuVmChMSuiSE0Y17vKN5FU6S/KYzDW2A6W/5O3f3jYwVg
CzrWq4zNnFnIzePhvStbicCBBW0hyQdejlukwqNaLHvhlD/Wnz3qq4R24Dzysdfh
wyaDyAtdcW/3U63MhzRdIlgfLk0MPgaQYkdnWl3Y/qGqsFZq2VRcLpcAtyvTkIFL
WGLpjkuQrkxQS3LU6WhFFXZqrkcuaLMpsaH6fhgo72iqCOuvi/4Wv76JigJSlRAV
QkPJ0tCJFqEUhEoMq3w8K/F+pLGs7jh6gewYoYaPNbjVgPB7b5gauOFlyx1dOCtD
afBsA8sufg0Bzpur32U5Tgyif0IL89sk7xx3eQCS4e+NxvqGpfksHYn3WFgd84GK
i//9SfKCFUIS9jkoHGSMKwRtQMuI/q+uAeebS8HuZ5yp6AbaQZu+fQbqdzGEFXYt
pYIlFS/2NHpsv6nJ0nZC+Fkc3i1KOXDZR4tqL+rkeE6jJz2x+zcXVm9LHDv0m62L
j51VXBM4zfZWkM0zswLQyWmnNAkFsWHHR43u2U6135o1RzIkQXhOf84kOGaKnkMJ
BYhvIbPlRq+YqilQi7ZycGT+R5j7UJvpYOCjCzrI/j/5axs95rPwcnwP8VWFnu5u
0ypqEdC/GS4Jb6jL7fAsCwykmVBDDOr91+h492G1esN2D8ogayw2fKp0Ve5ugAUl
rDDaJVw1QS7NPsJw/vEISUs48e2FfgcFV5SdElZakGD4mZ+R0vFRTPcibtjN/GRb
hy77m5UZ1TDGb6xnOPqT6IBpmV5PSbI+y3JGSydiDpBtERcfVSMN1nkA5EH6yKX5
3AtwQanHcPeITnhw8EawPL+OPs7wZqzqbYajGcIUlNdKQ8p2u4uRP4ANtIhIiAzJ
fM1yjhrBud17JHYiqpIyyK4V9T86vP1Ayv6HIJxcGXaxfGx76XwQZ0bLnOmKlSFT
cN4q5jzv07fBJIuQiekvpWEZHKg2/uIKgm8hzOjIyjhpbmBb/rj5lW2Qhd4M0zli
4JC5198YiRbYIjgHU1wuccW98L3BS4opFKD3/JR/Ffgw9YTTa8jGyI4ATjeyUWZP
a/t3yhcV1aRp16lsYfbPYE3YIikJG7hrNF/m+NZcqHPvtmpK2SnEO1DkWBtpAKM0
1T4WsUD1yRElYiQruISdNGIqqVoxZsHhpgHVep5+zZjNjmkW/oNU69wTO9Ij1xHt
HKC6HVlO/r/o0c0TzXe0aEE4T4Gd/h+O0Zcp2nKbWG4cH1E3xsdA2EUXnh5c8Bks
clDlQxMix9iBbpOv3PswyCEmxhmAd62pSbB249o1bZums37vI+lRaUsBK7JpJjiY
aZMXRsS6PauOTELjDCDy9b091waiHNUeklLVeqV+gTgEucwvrIo5JN6mrOZeBldz
mGDaXsesB8R/G8Du4oEyed+nzC8Z3vCJVLbXOwJ/+k03+ZPYfL9K7KzS8j1ldmsl
HSVWd+edYyjsZYWd/FarXm13ExJNLZlI/BCYkBVq+/c7rYkq/AtsckvczE7Tb/C6
VnxbvcxzZw/Z7rG/U2/N6eZG7pQeYtIynhpJxmsyh1FNRcCXOR+B3LDjo68M27op
cvzc1qw/uvJZcxkkY43xDEQaYfYQh7WQ6I9Y8oQTJqdIvHzuqVEsz2Nz3qCi3Oal
EygrpcUfVgTcXJxxCZz5Yb1a5JxX1cm0aroD7jQkR5H4G6BNhu+N9PrDRMF2BCWR
yTFAggI3cSqQJX601wXve/mqfwLtIBac71ICM9Ffk+OPNjTHBRqfwZoFL20klq7i
KhZlra9zs0G/be3OgEIJxu5mTGWh7hFEG1FJ23JOCPkW2SMNQtC9Ipc/N1GSLFqw
ZVVwkDvKl0XSOTumejC3TrVsmtppoytEjde4KxKIJe8DyS660U+zwl5DIKabiUaW
O2rjh9z+zKJx/hmzAK2TNR008Fj2tBhhbCg1PYa/ZZqBKWKvM5mCc08ZbA4bKwPZ
FEAYFN31Ik7aFCuo5Inc8/MlSGVTDoufxyvAziZwC0K6kkQ1a534w6ekEAO+01IY
PQShe/uUzIZj4GtQsMOrrJgJt1CeovMT23M3hxzqgDnBp11PoHhMT7zUTUuf8jlW
b3WgGb20QqUf15fAZi8q2XlOQXCo9FLPBFDYQL7dQ7eaOjCEmB1PTUIlrsKroHk5
wxzGbY83wizeD8plmFARw5bEtYo61s/E693d3r+i3mrmqs123OxeMgtg6xJAuJz4
VTSedm63GuP7ktW+U9OXZ2i5BkMG6bVq3nwBzcwNsSgTQlouBkzelrdwQb8i1X5j
IcuD6F4l1PG9ntqc6VVr3XKSBJ1ZlBzN+zP0MQLIgUfL0xQ5H4DM2pKqHTN5BVbr
ktYBDkYCmurkebskP8dW8GGCKJsXclAv8+1FMCqYmDKRPUjj66fYhzhrymqLdpqm
LMCMSc+hM3wF7CsPf7cA7pz6IIoULM4xWkhvnTuyyRLRNZYp8UppVLF+OSij2uYZ
l80VGYCAv7M0X4d3IgBannjoCkBiDp07kUA/6y61O+rYT4gSlRai4nWa/91IeZJE
TPZBkVd4O2MH90d+dquI9a4TZm0lss+SOKX8NuBYDJNfUTZcJpD6DDzPiS92wist
pLn1iuvsHZTnnSQpmby7cG3e3/nge8N8iQmXtz5oyVq3/tYexefv0RAPYqPuJ1qy
2kQW11m80W2BbYrvyaC44RfcSxLaHpWOCF8V00U6+JjcPLHR5qB9n1xcNjn+IEhZ
RWd7wRzxlgSpyvjRv+Uk7EWqVWxP+mA0KewD2cFin7N3NejsYqTZw+zpk/7J7BDw
6J5AyWQgSp5fH2gYTiZk8ICNk5/+wuU8tffzRLUrjF3De50sRvC0YA2ybCHpomb3
VoMuSvOr3u869BQeYR97VWziwgt35SBj7z5IGnTSNp7tJq86wcz0qDjF97Fiivdi
+Z76OJZgKd/yhv0t8OL5C75Msj7wbA4XinYUHRRxylDGBwZQKtktuHgzxSeRblSk
wCrqfEofMXKqQhwYyeIGCrw98YsD9tbVsaNsVwo00j5kcQHwoFVCYpAkXjl5MQDO
GMdONSEpyAFOZ/FJhZFkfg30FdWcv8Yu7fCV/+zZkW5eLRfIXIuKUpwMnIckqGOo
qfYeX2B+zAqGrhYV32TGx+KLMSkHDTcf43K8aexwSlURRERFWtEkEb7S2Id2KSUp
7hjnAjRtpWVahXVQJ7vexbQwXZ+llK/VkWDXC8h5/v5A696LrOEijlOYs1Kk6Kdt
fHdBTEGdvV9QPK7oe1e6islhFbGoCCmL2zXhU7hNXgCD+tkHQTmskI4aMlxYI+mQ
TWC/LCM80IQqLfHVx44f7uukHT3vfZIe5XTdjdzr4UAetF+BLXNXmc9hzMiADyVp
K3Tpn40V0q+yxwcK1cc4mdJLKtRRzgqaVjvviqSiqBkF7oX5nyM3QiIvE09HgBR7
zpgEmZCvxdxZ1NZ9/rzkwYhg1DSHROX4ylJ4rq79B6e/0ZqkpLuKgR0AX9mP/FDM
cSq2bBjY6xSRDvkAmjLK3zV3TpR/6I5yAecDaYIl/iR5eIisqrX75/xhC1ftlYgg
zYypkTHb2PSvEq2cAO/CTpWcZE+8SLvKsR+lYpoxbChjZjAsP2C7y/gt2x9xn/tL
0KAjdGIHk6CbOXwb+iGKRLAwOfAVXJwTM+GXXqsmada8eLeCERqtRXpYleFkhD8p
4NiXUoo278857TBW5+Zpmgt4seSCD+sP++tj1WuRiTgs/9BTp5hS8rQx/B/X3KPA
DBL4HGFhPqr8TknzEDQb+uW0SXMr/ygRWl3NmSXmhmpF1PzFm+zr2Em4wpPb7gYQ
NIbkRlIb8sZCYpmZ930LtPcD1ybmMHT1iDps7VbcgEv4FUBSG+3ZshOhDbz6MS3t
rS0xA7mk/Zq6XoJeswVx95dx1kGtlABEwdrRbWZP7d5huTbO6574/qAmHXycmU/D
jbe5lCxPc1UTHV+y1D2S6Bgir2bUogKb6wHHj2YhKYmOUw0my4d68EXX+yt6PT/t
488aAOUUughfAz2ajhFugBuQrjUp41ZHXMsnleglY+4BlqcHIIbVysBcQ0d7Fjp3
lH/EUCJlz2iR7NGoGdaUemqQnW1Ialk7hGgTI/7OVSjp8pqlwwGN6BKt1PhLnk5D
UsjXqdCZytBiUPrPAonSrto1LOHESroK1isAQh1Z7mHt8wa9Oea7hA1TcmiKFHwM
8G6x8crsK4DOjeVrwB23rof26pW0ErHIfiDtysWCiKYovO31jE5vz8Jqzhkvetoj
Jyz/A3gDsrXpJzGqs9obw/kNQne/ZFi+5MTP+ixysnZorwV+j+AHQNY2UonDGVlt
Kp0OI60N2EKmZNwlRxno3EQz1I60hrZfnJk9sX5V/yxZlPa6cvUrpXtGHF7/4KND
xKNlqtf6bOEUJNFUH8MRtQJAWfSU2HFJAjxRjI2KGLcmD1BtBv8j6d7x9IVwTume
TQlSr/9flCde/avHbPmIhWMS7MAoz/yDeDIPFbuBbUs2LMMF8aCluTmsT/HyKuRx
2ViNTfD90GcgUvXAJEa6Wk+WxAriEOBzVQjOyzfwNR+p1l/uxnzF4TngYR95oyfH
nCp26UTh7Nh5DwhHsgHz/vf7yaAt+opILuvFpXAMUmK2ShgrVC2xXUQdVl+V5exi
SWIOR4njYB8Eb3FrtSKqVHdmx3lId5kZiVS5WoTQK6RfiAnBLXr7o0KXHcQ6vJEJ
4nkrgSvBNKXfjure5pR2dzbZ2Smx6qQ+rbPh2p7zFFXkoKPwMPrAwt1MpogQa4iZ
9CBm91WBKKvRxZFbdHkIKFTy3hzjkSDFrEns2hhMHUrCjfKQcNqb3LLjcps+iC+A
IwClbhAEnXX+jxFGDXRiw861Qws5A074jOD0TOcczM8Ihn2POkdvCoG1WJGWxwHU
z6XOjSu/Vxnnte9902TCwK8ramXu7zz9S7PPQhzIxzVG+0eFfNzsxCU33wPvTa6U
6IP4HtsrLCA9TBk85fENI0D8TuiQsg1tMv1QGDkeTk0ybj5NxxK+wSPlv2ZLQ0tg
p7eyDSM24MjFfYiRYQHRag2VTG62dtuaYhFs6J8VRpwHVcKA5MG1CNtmEUqp3ZTm
rAvYQD16AkJnXtdr9OkYJ8+jaocA8MOTD/tNi5kbWH+yvljT/COQ5k+5w/6g7gic
2ktJU3oNPKe/vnTClBhSPgoXjdBEYJmLHWnHoPlbHfYPqzcfqXccYbfpviQlfDGW
DmsW9jaRydmgz9X/N5xOkMcS4nMnoUdaP+R0cWQ0FSyei/XTSqyZo8CVTflG7BDi
j6BWju08aTUssvsY7nqDauQEwQA1lxs8kzJrHegKnKTk00qvXNrg8Gj2+nJtMnwH
5i+ngdaGzFcYG2h2MjzHP2RhmCMA8HhuPt0tROngzF0HMAZwoOP3FvS/O95jYxf7
65tHU5hE9x8FYyqgp3SHcy3LMjIfM0wiiUp0OJPOk4LuStLlf7XVuGi4r9ztUn93
/l53akrRqR2Uw4+0LcF1u8hc/jNBGkwZZj7k59zRILybd6JNJ1K0PYOkvgISXEBd
Hqid57dMm50hK3YKvSFRBKs3ZTmPQ0CAQ5kSjNFHLTCwKAouK2QAzYRGmQXyh7d2
aeliJCLFThYKz2ZcvT9HpJHDxclku8HR7e+/wXfthh5OLysQZzrOyu2ZN5B1Bg7+
u9PIJRnMLZpAzjjENDC99YSq3nflP4QM0VTP07Df2qgdNNhCbPVS8VJ66yb4tehI
ULr6aM8tzdX7q3/MoBSZGo/AbV1pv6LuwtIFAwqDYla7mVWGNGzqkJ/DZJAlfWcE
brqXYRh6Uxc2sJXkJr3HV0ZDdYYgoXMZXPWZtOxTULf2bpp+YN/TBTh9/F6STXvA
7aQNOfdV2wCSKYU+YzSh3Vt1I448lvE9xkKxK5xi6cImipaHlKiiejiUXsfBAYTC
vSHfiFbWk3ytwoeBXmPTktNuwh/eA6DFaysw/s9wntOlLcrumONSzJftRJGNNKbK
Faxwi7vB6+rT4SKh7e9tD3AeAdUILlrYmDZFfeefKfNvz+YnIv0+WFAawYZBku50
HJAsU8X2FvKTPcG/oBjcSib1octSIOiRRgqEe/ipi1wAse8mlqDmbF4zAl1WR4uu
o3j5+41NTchVLJuR2Du2Jm5xhSYCHE5fchhVx2ja3rR/BdDcEoZOEKKEtd31G/nJ
t8tNyBqWGRvjOOi0PH/auZqxPlKz+Abxod01YmJdrCfQUEBCEf7zYFHvWQ1+B5MC
Cra6cly113ImO3+P9YXSErsMSBo00cscMxA23Bp9qO7y/ah/wicP/A6HRdmv2EXU
IfTdWcny/775Jf9RkiKU9czIuHGIjjitI1Y3uhdGXeObDxyLbPJhD89mRSrtC7KF
mqPYhayEQHd6aOee1L12VToFejOo/kMjBtAhQFN5kjU6Of3Xv4WBinNUiMdafL7T
ubowThnAiOPBNqSPHr7NRf4zWAPgpEiu6gQoy7dU4B1giZIBEauH54JPVcezskzV
EFc6CHbckKkITlHjBYlitq1emElLyN5UcGI/wKFsyfY7iHeBhwjBmOLdHLD+Cikq
hRcDMlf102y4ZCkom+pOHSWhjqbSubH3VLWZ9RwMNLT/EUatrhC7ztbrO2F+i/1U
tZR7KA1uGN/YDQOKpOzqbSBp6lWypaygyNG13IRjtt1OmBH6OnvYYNrU87Oj3tKg
4orjUC2URR28RPikDchAW6Kz+ZxrJRmTnXArSPqlEEHOJjUMeNHSf6nHLd4n1XQF
1V5N5dxs7TTJi3e51CQL372EEcsqjXX0dz52erVPet7tyeVvN/oEBcKJ0sAOTZfw
ue6sk2Epmr+AgNS92PmzVx7CKNFLeeauTczev9tJbLn2i7xwDFl0PSbJ9wMUBy0L
lcC97DxVjhg9lWAetg4oWXMh76ehdn354N33oKO1Ja+mLde47tGk7G0uUNtmfO5M
cJdpIJiuJ3CoKLe4G/3NfPC6OlN7I3L1DUXPXmYgjbESskbrB59JD9divBmIekbY
6koEGrNmO963qZzMOCgvUIDlrnOcF7tmvN5su0Ui+u//QApvHedEye7z4Tg4X7dJ
ARv/Phst/qqU1at1gr7TQvoF05iYpJiaI1BobhbZ78UPifehGOZQePW8JExc6QXJ
jTJq/36V3IVwmcY4UXXJlBzcetxZEgpUDhbufiKhfVGaI8S6LhNcumVkD+d7S3nW
R4Ec6IBgTuXZjL37P1Ce4PDQwMTn2XqJ3Ky1viFnnTjeYhGWN9GIuAG5ge44z0PZ
ZzzPm0s7xya+Tx/X7meGtz5tJf6yf21AfjJ5imJPPr8UbgZnZhsuXbj1RwbYPfON
+eAI9n3rN12b3NVv8Mac2RtoXPMwn8u3TWkPiIyV0fDO7badq2ZOSSdi2CR8mdGM
NCQQmMcN1QTi1kIt4c21yL+Y9BF7JI7LAay8CXzmDUGEw1kkYdvw2l+qnd7Lvhwz
hy5EsWg9NBZ0DbyhDOesLaO0z5lkKnVdNCfpIDGje8p0/w8aYgsaoElNva4Jmdj1
SDJMGQJOUZRrlINP8zas/ZlxRpAu6HGNRRf7T6aXnRNRrDM/AVdzET6F7YhXUbky
tOS9vRaWgOsey3Mm4rccnGrwLtYvsv6rtnp75HrXsMVmIzYKpyiAa2uUBkD0fjjC
x/9RQV6U2fGtN7LwRY7JBUgnu1sMOE4eT+VnLHf6sikTno6iDFngKGq1lpne0CcL
oWoM+OCYuV/BlQ+Xia+aIv492iIdwWrCr+rQwN62UN6rIWhcRXk4kHkSECyyI3xm
3PxqmEQg+d947MZtIu8wZtwmT+lshzw4A9lEbGWWxdGHCdw4P8VbL+cDMzK0sdfT
oAYHZxTz+kfm3bA1+ucZpJvFPZ+pvMLsf5d9jk9j9KEBNWbKdvNTQmgXOZoBfuWu
CViOsZBvaj4XCD3RhCM7vjiGA/YW6PPJ5ojP33KPTpea3HK2SDAoJNAir6+TU24T
ZEl9UrDJEN9bJ+UdBfBjnssbRBpKSA3ccqrRnuqmaheul7utXn6dqiPuhuJcr1Yc
WovUtqdAvJFvNA7MSKqVVRuPCpbMwEQ3sV5yCQNRI1ySL7GMp7kjZIjOCyePMnRw
4ieu+RP3oicT6X/8A/vnwsEloQ/kTBjbtLy8CMBAU1MQ/o3qI8wYD80yNV8v+ScG
cYS36syxb+4HqVaxTB2qI4RHVG9k9JfL1CCtGLq38RZJKTRI4zA3QBzhLRa1wZqx
GESG12rzHtMz/Rl0F14EvQf5kgDoiqsnkANEvE68aeIFyuWgkKFgwIt+PSnojNsY
8hUkCpZYUbGDFo/JyG8+HqM/KJh+HStERUe0oz7rnnixCyVA7W2KaJ4rRVRO29XH
ZXG6L/9vVeoJ9WR4VEL9vuF3Q9lp6h4ynIa5v7ybVU5tCP3h54sOwZ4mQ3ejk7jA
SlvJ1+qXmjZgeWX+BV1nqYUL0vY74bCcNSPACHaI6BTIEmP9bK3eKjeHCvp/sA8X
llMzCxejtrHT1jEGA5WfklsUzbDTtPU8tu5Ub5hPd7lBc7ZFb14/tDl0z/avkLDg
jzGaUXns67F0qQJlXCKq+qVLOv11LJgn27CRJp3z4ur+6+8qmyIlv0NoZu4D5Qmg
rEIr73hB8grf5ycEry7SeHRYUqiIGlSh7wCgOWKsyKml2txfSBUsjH/wyqeI/AOT
if0g240UgTNxwAvPiRcO0c/BHA+SOSWb/xBApJ+4LMg+OA8C1zu8A+CbTxuZROqN
0GSVcyU/jh8tFu7s/F30cd2LUzpWcVEH7YWCwLJtJE9xkxd472xvbVPVsb/Fun0B
fIpmd8DOFXtLXJn3XMI5eXT3bpyEx6KZYajNPxyF5uDwjZGRPH0l0UDu6I/cfx7W
cPxpNjZfuRNJvMCwnnWWr0e6nVK4FYuG9u4eBYxPiSi/2FTr7s9Vlg5y5S03ocoz
jC0v0+q9oK3q9NtJVjkIgURicaoIS4RLUoX+ZMYBlnEjHwxIN1V0OA2VBGRopl0T
sUrk3zeltj2yG3zXOdw+IPGvxVEM1mGfadAy+Id0/dn27ePf/u+J9/51kr127FFd
MOCDwYkCHCi/N35YpUuLyEGqpvw6nXxTVNHORhoi7Jhyt0tZkq+HxRa5Sd0c6rFj
ziZJ2Pr0ApHm6D8ods1JQa10ZtAngH5+syGnb9KnBsCBMIjZ7yCMPo1ovVx+PQpY
ZecEPGHh7pxuhsOjrBxj3PGIUarQcKO5CFH6aL4uOG8N/+u8Ftx0a6Ct+MNXmamz
QXsrmTGR9VdCFEzzgzse9MKYS1z2FvKjS2K6tvjn1+kme6XA+EDRlQ4U6fZJEYf2
lENuqe7qaav/Msy2aoBGBt4sdatx5Z8yT41b7kEC0W/bhS6KrlJpDUsfNFdOquyw
X1hmOuyC0pk38g2yQ2RIx2jEi4p2hhx9Th+opoRYqciTQ1bLpkYyGZmnWk5RU4gQ
48VbbO8+tqqZm0wURKqGnTpYcwB9spicCThNvRCbnNLod+YRby/fRJ4lvuxYPVrY
sACakI7RuPtNVNNde5iVsrxKkrAhSeYmS4TuoJAzMOdEOn/+cBuhWs6T9Gx3MAGQ
QaVaRlz1t/943Uky0R2zCeSC2wFSpsBU/LBrgWLCHTUaRAbnFtffeMQGRt6c4Y9W
idI0sqZtODZp6ZEXsi0U9DQ3lRZrgtNSlesEIa/I7QpvDEMO78tcl079/f+xlwbw
La3pyVzwEsUfEWtMVCa62HHioEOEb8vaGaLh7B1/mzWyebs+cKsT71grn5KNtqnp
HI+oa20/FsWF2+gE1Q++io1U4nVYPaWL8S8oAeyPyPLjJqEshHwsBOLoVbXO+MQS
E2Nt1OoztHogd2SmwNrAyCnvp2r2Nq7hss0tzNEPocwbu0ezg/Dmzm3Fo8MHbNaK
KdqrZfcur8sOQ3XTCUMzfEK9N4JQPlD0wdNCxbN0Jebf4t7RRTovazZ6zOOQ6pjz
Z3PBYODya+OD2c7r7sC0leUAtMyEu+MDopsV0AVAO37ymikUFGepDoj8QCQUKGMV
XYWb66E2WyS1T2sXWE3Ml1ceVC/363pAIJ1vv3v945z8Rk1uM+IItC38IG3KL2AN
eOtlKsVSX6qt0FNBbCX9frfhlUoiyazXKJ5VgPCb0TvzIiVMXchoWI8m2KG3PuTy
55EiVKaYqydUnoS5hOJu6FefLq3ZoaXWUbSRQRJrBb8y63RlOl46sQBWViXW/p05
TphAbbhZWqREX14U0soSS/PsQMDG9uxkY2/EVk45WC4x4P1VT97cpue2USYjEFJz
FC3C/zYmFgnoHKOa0x5YlrDF3jOT4GYMEeLxzov+Tw4V4+8Sewrkc54SZHPrTKSx
4TMMC3bFNFHjAC+f0cGOrWH4CWu4FtjAbx019iR43HirPNHOz4j/3eO0Ao7nSc82
tUu/FABdlMHpVvX2WtnkJ3/9sVb3H8Qc34roNLNfNU/ql4Ub3OLz+2XzG6wLOUnd
lRJD7++XM0fpuePqQ1XvMkIVpu/TAQGgCDh3w/GchqvRDvmpuPxPYL42hDeRIJs/
WCiaaXHeEQ6YEh2ZpybkVpi7wJkYXstDSReAz/aNqiEm1s+7WYEMrTp+NpvodToG
FuMEqpDPAVGUTUBJ9E8rEPyE8vuOSbirs2YN2rutv3KFBoZyJny4jbbbagEZS97s
IowQhAe7sc7iOrjSnzjDgXITnAQZPdNEccUb4WA/VFQQ24103Adag3K0x5It899z
pct05HhYotzsv1gaTJeziTRU9wX/8VwcGrzAkQPQClRF/ADNHVrbHz9Y6F1dsTaT
oBw+tJ96SZd6EACiifqmnj1sMcaZGKwLZrS0R57pXSWnSNah6Gj2lQryjpogE01E
klc25XZGi3pvfdmbrIkGgV2ypy7QIj9Osum3xSywvLmr57/YJ/Npx71cv4+/gvgK
PpiRxCA7tvcykRcN9qqOiJ9d331iyIKOr7Syast/hb7yONNXR7vapWZY6m4oFUDs
jpGYxBP/hq7SKtPjflG2YuVyc30lccPjvWnqIc6gW3AvqYulTUXl4MdJMX721BVw
A48NDUaIDKdxKUJcxHE8yTTGF5A5Rwr5MAbl37BTdW61zfvJ1SkRd/TYGhAPOcfz
ip/Av0zNHsj5BBPb4WNSkIjimzHwEt3Yn+jUo+cME8e4+MxRj8GSlRnEtblyBOEg
XOTqRzvHMAFlmv2BAm657VwW2HS83k4jtPeSo1LG9jERf1hxmJdaZwun9yHWz5ut
e7ko7mtrk30WtHWPYnpOaaxQdRy7fJObQU+Phs5PLVQ1n0KTRUHrNBbszc13jZ2W
jP1BAu+7JMpY0DvjZv5I+7b3q8deGktPAsSudbl3AZLW+ccShx3ynuBXpl+XMOFZ
l6ApcqlVApz/6nGiXgBR9osH/spdXtJ4dt2HqOBS9rzaPTBrQE09gL+o5R1orPnl
5xHWQi9h5Js21WyXs+3cxqSWO0WfGVAIn2EWixoTJEQaGAvvVW+F7INNX7qFSv8A
h1mjTTY+gouy0ST8BaihQzhsDz9/JKVc44WEx76XOmSvC6zAUannDsBZQiS/Ut5G
gIBar41evVe3OZ7pPNRaav+2mpRu2+iiKrRvuzvTg6vRvOz/DWR272X+rIY+qN+W
OpVYVqnp6yHjhf9TqNx9DDBIXJp+W+u2+VPT5sYjPI8aBNyfAATRA5+WUFesPu87
nkqge6VAXKpwUTVHVVZGfJWOfGoAKrZDbvj4mBVI5lMChCQjaOuIuqDK2Zugu21Z
Iv0A+O2wYWjyUgwEXH7GUuPjYisPMGEDRYjMCex1NP9m4MRLZhk41TmpBDj/D+Ul
4X3VHf2FOaRtA4EoUYrnJqyQgbcJUYK7gQN700SKJdXf8y/VDzf2ttCIMPZTEgDP
S4GPzAQ+BP3SZ7HwdmnyavRGPcoraq3MDohL7ES/RFSd2cgg6geTnngSXI5F7m7D
iryAXxxptXxiCgTiMzT4RlgfYNr8yko9ime/hXzVc+yO4OGy5GCKozBX+RTAwiTJ
eSbYbUC+QQpDUo7yCWUo1wWk1997QvmpHm+AVZ1H8OePJxXGKSf/zpgLEURrO+8A
z7lsiMGypx0XtVtW4MMs0BbUSfkfFnKLJ8ZKowxt6l67mQzTEP5Drd98u/pO06bQ
nVnNHjJP94PfD+i6Cgdwg8KQqqSROjrPu5CynFYPQr3YaCXesarjjSPJI+AanuxH
SabaP9cFl/tJfKM8JSZzuFREJCDikg4IlQfvbSC6ekPXhNUPa+lPtZYLdg6j4OEQ
mGFFLPRpfkyU8ShFzg1sy9DZG3ogQfjdYEJvzVAYthHAdt0jTqdnhUViacCkFkY3
zFit+YxcYc00ObngxVABbAI24VvQ6aVQunEsIcvvFfOx81XE+crEWRbdqVizzT+7
GhJ2jQnuDL2WqK518pRn3kzF9UXDFwgXG5BbjcZwM8eQhoZqHjlL+I8e9KKE98SF
sEz05+Y3LidYgaKP0hrM5/NE6/+xN+5cf4uYEgR1UtP8vQeKYM/BUBCb0LKr7R3d
EYf3WqBvTyjupPCxAS0DhbupJ7oQqQ30fyOQTjjGQTTrfb+1LAXAoIKGYMK9l0mX
c/v+pIRLYeJvwPUqUF28rC3AD7Jkus+W8GBgAoPC3fjB8AYlSxBxSrH7eHhp/a9l
ois4vDAmJYpU/AF6PMlMaf8aU6YXbQ+8zlxTWGSUgIv3uK8fElIjumYm9ofO1dUC
KGlpjqZrUnnXOqUKbB4PaBx/TVJpGuAIKjlUufgu99g2CcdqZ6xUNemCP8YSAAMd
OR0WY9Vh+Az2UF7iiEOatTKWLWy7+FOjUYRvAJXG+fJMcEKV4KH8yM3mLY651kXD
YoZf086erL0jMiq1ME5QnXksGDTswZ/ruWh56VuwO0oGVUjwfVcruL0WD0PF8GJT
sdC3zftBMUfmYNKYkUUBo2/tWYBJOUs+RwSrRgPSHt//FkqN+h1l8wcPOAX2E8zw
y5bkWWhZZF23XDIpdknzncihY1I3MGwvyCSZobxarr2SHLWq3gGW9maaRf6XF855
wpui2NoYuEK/v0hhnkEtVUAfnnPd8jQ6YJaePQF5o71G9jaCytV6+pNBQ0VJ2muX
Vc5VIyBeYsPUMPBjhbaVHRUkFr3npMNVkICrsO+YUbIs3YtRN1jePRABKpDB8hY0
n2dpWjhwB3kG/4XDj5n7qHNSK13LaDm8kU7vQAJnH/cUhF3TUAn3I5TGgfMRNw4U
7Nz15DT0aEp7vJPq7t+ooiRmx945RoMs9r3HVciJkewUCjGgmXIZgx8uJwy2kRBQ
5Ar7IriEinEBR0nzW4Zw5B6mqOdKRbsWdgYEauJbUvcBoeDkGRQmWYcHvmp29VNB
UrgbIQJmbGuMFnEU8M+EvD6RffpcE8PHvyemcEj+T9iDJT7DBeUEU9tjSIWnjk9f
55pttymdPuKKYAZ0apKdu4keO/Kf8lIvkYIJU8sHj/vtatnRRgq2ISbQs1iBYtFk
y6F488mnlrxzM10E3c42APIZmSpkXmOKPU/arxd9wO0Hrc8YCRzWDVxUhg5DH0En
Z20FkgyZSTUTn3/a1a9tiMOZ6UlG7X3jFy9+dJA6pmyTMCNH4LXkOGKNsrDRaT2v
nkl/EEtBGjIMXPPS0rtDSGvDaIpBUSTLNbZ1+elAaIWDreYt1ikkB65f17k5MUNX
pc9KTejYPRPq3v1n6WFfu89VhgTlM5Ge4T5Tr1EMnSH66xDWWR9BA7vZrfk5Oznj
AZsIn0gEtH0Uyzu3aXkkpxoBeC63YLFKpAOvn5e2xJgrRTGptTiHRkj4dvJb5Jep
2ZmbTEsiQByl6Fapu57vHKLD8E2LDaNx/j+VFoJmuZcByf9UDW6yL6hRDxBlo0Q9
t+G30b9KiZNc/tDq543eeOUb+4k6tjAFgg+DBjgzOzL8gUUy9h+YVUrk+nHMqFu2
+2gqiUXTdSfg23Yn7suTJ9uI7S4Z4BAEFYLdrwRPvGfsenFYFATyNTRQrOcpG1B1
RlNaE5BbFJSclZQnNDNhKqFCdGIb6KsfXxtgYJNxPR+Inoq5Gyu/P86I8oc74OuC
gUe9qOzWHY3Ks1vbUIAHQwk4sP1p24Yj+q+bDhzNeckGfK9NrsyuNRWsDBQUhFPQ
vAmTotj5WfuwbgaFJONyrgTj8xMWPTU+EWij03QIG2zXN+WeeHYXAneWwnXUcRBg
rGruzJgQy1k0PhA8J1cexX6iX6B59uq8lf8pIf++L/6hUSAkY12MCuKCT/Fq7TeV
oZv62pVyMpy27fh1Bwj5x90Dt6F7QIy8in2fqE+JU0TRnntzIJTUQawudhRjkAyp
DyBx+uVBSrX32Bic1TPWuxriY+9m/fKBqXmg93AydmzwuXsK35BoNlN6SlNsfLNg
zvlE/8Q/ZEP04hELVgMOpT0hfSKoNbcgp4uFGqU5l0OsciGOdWPsKT6ezeuVicMD
y+xPUeBtRutSTxsVEkYhbdD9ONHxnVdxPInwyrIf72EyfMIUXvVOJHSPjp5LH+5J
Qm5Ypy9ZfCvgVR8XzPqO8xk76q6FOxXqESGYTj0ys0GBH5reKTFt7NO1JNMX8EOP
1+kl0vrROHcXQBscMYGqHatfeqCmLSTUBdY1ujcVGC9TfBeQ6oRsEnG98q3Xk6qK
AGnjQVyhvcDj1oKEfa/mmF4YUegH2keR0JRJ+apbf/kLugCaV32qSuILfhMki7AV
hx4oK9UoZpzXrHf+sGkNZqWu62UI9FECM4YPIVK8RJGDx3MN+5zmanwkS10yRb9z
7ZJ1Aep/0xFYJugEfd0l3p+dHYiaAMYeL2aoQHFjKX9Jt/oQDpAiuNoGHacIePLv
YEmsFUv6//1QYd+XzJGg1z5vO3X51CmVynM4QrG01dvF1vcQ//Mds/2a/ITLyoTx
fxRkF29T/cUIgkJdlzdz13OmHn7r9MHlCwzBwP/Xhqw+3svWdqKVDTbP3kaDsD/x
jRGsI8wMLhpUftmYHwcF7u2rVDMEfygyZBhoCUlQvlkzIQi4shCr3Sc5C97XIRmJ
zfpDEUL6wvo+YNH9PzsoVsT1lwtfgP2fa/6nKDTe7lvlfmilgbaa2DtJeLLVmoHa
UEp1YzdyiIKoy+yGZnNsOpsSlbpWZ+FOrmt44y9QQhLyPcogN1Mr01dWeMRJCNmV
7XwJ/vy3qYl38DE+3bAu9dar8pooUSwSKE/wQxRe6hEJ+eSUnD4A2bzbvBY7AUap
v6MxgLj2pHNaRhCLO1zldinAa2AV+MIfazj11ZqzutwMPEMCJQkV6vt7fVfC4r65
yMb0A8Rnibn7FXOfVSIS03jqmrLZTLju0t9ylwXPAE0TmlfU+7bD4kzSvdvWkUZV
Pns1GZEWcqVMn3AwsERD396J12pcwK53zK29/hRh5H4zrVyoA6czKuvoAumdwhNj
jlKOOWLiDpR8JcvmF6omsCsCNZEAn/T1z6yQ2LJ67OANJOz2enOEFezzat5dantR
1Baw0wwqDXpP7ldTP4UFTwz1zO+YcoJEg6aVx3kv27LvOhvVwl7Ez8hbtAiVzLAU
+Q9Cu81hMYVACPBlqLf+6WeXG6Uo3UX5PINvhvenqWWPi1+GYnle+og3vbSB5c5l
g60HC+CGg0sovf5vaS7OVP3tKk/AXlnECQP5uK5t9x7n3kipz4yXr5cbejcqcUJA
dLLZTs1gQV5d0w5vKvbsA0SLvTdgx2uVvwNDJMVDZ9NdWa7hRa/m7MPosFx7Wb57
0TgGvuTIGdNUNPBqszJ2u2z57uXWX8w7CdPtYFXcJGhJdCe0yWex7CTGMnvTBhaQ
7nPTD4QYpCxdVFCY3HGqp2Z+EeF8zC+leO9MzrinuuldX7unbwhWOc/wZQ5tuRuu
cy7WjT27vHdRTPsOrkD0YMEFOcy+lQURH8qXgYBWxsXlAryQu9ePoO3JjvJg/6qM
0LBGKGe9SB2vVXEbsACIZBQw/USw7FL2w6c5seh1nr0mbRCwLYcIK4KQirdw/mvK
QL9YDTNhX3hnziOo8ZNkDC0A7IwGX/LQrR+a1hnLvMiz85SF49VLyKtu4OOWTAH8
bHs8XwnL2eggsjAnD/CJ4LDvvvRmY8riuqx0piCPvg5FEONoLLE2sCzMt2WNC4TL
KHTTxAo483/vfjj56t8rnQb4z17QoudybYY3xlTDczkJyNc7vFZqbGnMDw6gTvGY
LlIzNscSM/SnYJazZX4KECx+qidWSdUxLGrSUsHFRjZryk8SNiUEXgaceDzL2x9Q
Ak9MaOMJYdPBiDjIFJzdH3RdddR4xcRKeXjY83Xn5xBqAp8jaCxWB6WZDovJ7B/o
c7Hbz0YDSTlVcQeGj6IZnmzXMpoIlDMXEuxxVKNQna4OdRwEbaq8jHAJAcUqSlMc
RWOEZ+OTbcweVLbA5f+IPfW/kr34VJv164nJTN8CSOw3A5978kWXSoZgUBxJ0CN8
tOioLCFYybq8HMY/8GpUpFbH6zNJ/l6/iDrV2iA94ht9eAO/iNjKbV8GYQ7hIDS0
wJFVdQiUDu7y1uDpTRa8WuXhu0NX2ztN7lBCoa6jlgpbpBC11Y/666mAfJCmhgLl
zPbcUfjJfVXksGDdymJ4AcHBo6K3lud16YXecW+Iim8gcUDVwaKy7Wlly6DfPFPD
YgthYdA/kVTSaVcHaLMk8kgZY2V3o9QMypNKc6TWFB/kdxux9mTy/pplgN8Jgd7y
48m6p2Pa28gd0lJ8Omrq/GbwSsTBQu8A+xcvnmtpea5H/HwjTXYBwD2nkkchs2zS
9lk95W0R0D8whSKQAbYmmEF3uhqPzm141HFjrNm+Dvsvrf7zxReIuVySbL/QF5Ir
XAWXVKOjXAFjg2pgVa76nZKk9Guv1raSbpA9KypBfugyClmnf0luQRzkpLy9xZas
yGlZYrEako2P+ITy11EQ/ebnUV7nZJHAJqQFQbnC6sAE7ZK5qvjp8jAFhNb5GvPw
fEMPKFQHguEblKQ6kTAYYhgA1AODXXN9Ks5ch80fcevy+6dus6SIhAKiwBJ/YoAE
MqkWt/YxfhZDif1d5bG7iDyk+aJ7DubB2Yckred9Zya5wEyciFizy85zsCxpvl7A
zCKc4qbHVDcQ9ywpb1pLTQpkp91bzNv2UVdF9YkGzoVGRMnCMbhD4iQLMKI898DN
SHJ+Vh/AhL/Am6N1ugRQJ+LtS22A6XO10wrRC5ZTxzQXa7wkbKXft6Uf1Ki2qhb1
QUG7aHwODFFNybuTz/vrwmH0dCaOjKpRJQ/L8Xj/M2Ej+5Sg6rWoA1U4kzOoeE6s
wwhJ/b91ijRqndI7UzMct+AjvgfmVpTWHYwO8/gg+bW5zerftaCqh4Em57eOFmkZ
4Ah2ZR1nO070bgzqMhfi1yjDW//C3QsCojRMVcfdoEwBouN+DeZUqLChZHejLsOG
II78SWWxvAo3leNAw/fK8fmMOuKb5OG9j9ZT4i213RDnP3d0BsuDUH3LPouUbYGI
bn9KJt8LBwdwEZKwD6Zgq1b+hkZG2qkF8lVUKeMhs9FPLdPfe5e1mEbTjmVvkqqt
4oULirl5uPIorf/DgGRcnU6jZtMmasS54c2QOMqKGSF70eetdpNT53/V4m2T3D6T
2mtB6ftNGX1m+h9xqQhoI4QPd+T7XvBjS0HxsvOJfgF6TVJic7/qZqeug4q639Js
QQChPRUOB91kqgeXmb3okKKKQHaNI+VtCUp8r9u5ruX98USMLaOVsDweamXOQZMB
1ufplz8UbxFOLYwldgBOsWr5wl/hPBx3SbbjWFdnBJUhovKQ3P1bCFPqG7tU3Dla
0Ze+7qKV+S0ojZsBL6WlmoD1b/EtoDJLVHp16nWWMG0aq7WG1RpOAUkksoEvmKwM
mkcQn+kZgkuMLjcvXGOHgvMFqLVioM/4CB+RcF2xlfJhU51ACStXZAfCs5ELjzaX
3JcazramhHyA8ekOou2V9ezGEkABTppTsxM1jRYTHm20WdNgyj3WK5AunnP/bm/n
iLwfyGZD+yvN9uDJn6WYswNpnsrZndR410QbeUtPHi5s71/I0MDVbYR7L8gmrKn8
JMGUQbuZhqUH8Vu/Dvo6nK8ypycC7TDnsRNBKlh53xL7Xk5ToKOHA4O3GixB40Nt
TH4PlbHTMIzlC2WgxKl72c952R31wKykkRf9IIN9e8ddxwKEwj7qKIDdWD5u6xx8
4AfQKZlgBUNDNQE07BX8u6JqDQ7gVdWQClFYM8wY+FRGqutKqW+g+HM1VJXCc+NE
ByKWsWX8AVtBSuyTuqwA+1iI+S2ByyAhpLknz6HRgZyzfnEgfZQi9wBh0++5WR7w
Al7sEc/Cq3hAoAWIhaclISieldkSfWqzj9u49LR+8AN6Zf3Xr7xyI6iJMWKhzUlJ
/CjW8WHmSmlG7IzMzuDfjIZVnxghvYKVMJnIm8Gui/M9XpQsnkltmLG25HPfN8oF
c2WH+8ekIAvSp1QI2bKSwDpQeahpag+3OqUbcBATqMh0oYcN8s2tRWKcVVMKaX5G
0PaJyts9XGkZ0+FM3aIIlSw3irfeHtuSc+2/0uvmombT17e/f2fUYIx9do3Qn5kq
dph2WF0HVkZyQMP0Rid8sZVNfIy6sUEegeN518hDRcOuN2qelsGD+MXen9/N9jrg
BHRn4AkCRNRD0Mt7xmRgLUcANmnwiPb5hPGAsf/FnBbYF4ROvxRsrcEzwD3sNp28
mdf2RJDd+aliaY8hHVBQ5I0kOpheeZ17S1AAMITVY4blnxdDhbKIiOp1Jpf70PAK
KES64MHjRQd9jU1ne6sGZOJoaXV9wCM52mLQINYeQYnRh8iDLwRoG1PP9d3P38jA
S0gkk7Uy9aBaV+p6ZzFBsmxJoiQgGn5i8TorxzPjFrXx8tgH9JkkmcwQcla1LgpL
bIXN83wn69ox5LzK8o4ivHISag/Q80AW4iQkG9hnbJ9A8sk1joT6wQ8MoHOOsl/8
6GqS9GQCcAS/fCcVdLJ6Nhhfjsn6f7Zre0nGcY0i994QRzn9sRAJCfa7FTxi7JF0
lZVj6J9pkXWjS6+WXTuLfjViG+4KXU90rjVOnz2PvG9VHzBA5G7v8k54o4cyqOoI
9Fkb8etLesaMA6MjAO6Wi/+/2vmHDCdLDhoGgMh3HTFpdZE1z0q708mxmBMwHtFK
5KQiW5UQeEJXIIr+owim0DONDe9rQ3oasNjStVukVpg53RnsRK17VBAn9pqE70np
ajfc4lLuu0k3+2SHb6AA9sOlX+V2MGuEJH0FQ+hB8A5OMtrjdvWWJm0L0vB9GypN
ef6H83tGdQDSvbCNnE3HzzPJ0XrMaHXl6Qfc8g5QRs4odsGBilzZV98Z7MLxOIqI
DYryz223E9I58WhBWSsFsrP5dOWXJCPbv8KSWGFLxL4nUcXcJgtBGbA637nUzrsA
PO8YpN4Q//91ShjuaT6m9VXNxxiWKUfGiUec+S4l3AQWwDedkmhKFT0WOb5QN8cx
GWgb/JZU5GJWm3vIYN0PQSckW5jjBhJqOoBs2g+9wSBFsnjY0kS/z9XrFHxrZ26q
lAZLrM288g4ezcIw/xZXBgpd3UnvQdP0sgA5P7odPWc8Q2+ce+JedrfJz1pQCD5h
YwYqRtoSpILFCKaYWoK8amPCJ+UG1FFqpHG6YI9X5jpAK+NpxXwXrVysxavVXg1p
IEcFtS66YFLhcRlx5GE+g7AOIPCu6IStgXExY2mbyiWgXkI/05rWoNAr3sA1zyKL
op/TXl76LJWwx9Wu9ptoysTXBS+gKwtBO5Nmx+vUXN8PyEMJScshpswJq/yujroT
V5gmDleNKi9qK/gIJXze/TULQ+JiF+yGcsCg3u1n31rCD9SCLxTKcRx2cYsam+/f
FowydWcJ7nycM/ryOswXC0HwVYfddNl+RVZKAv3l44sq6i1opuy6QUdkXHpGttZ5
B+m+xtnULN2S7YxhQ8xh/BuNqe5D9jmi/N1e8B4M/PKS/aeiPL0vtH3xl1oyzyya
bJioUDQiQ+AfioKUNiFfy5A/umorq1brSTTeNaUbSgXUCrZV/Ur+Tb0Joj7JNqTL
/kCh3T83hxiJ+uAmFIWt4cRrGLuBbuIpbp1LQPonYy08hfejQPQ4+ZsLdjCg62Xi
f0xYVF4YRNFfI+39/xU/kNQHWEhvmXgooaPabOn6cinTpJGgXaBF36hAzJPQYQBA
ubQpQQsxKGEfEoRYVIYQnIQk/IcAec+WEZwdjapmuJr2OiT1pRbgX8N5CY0u/shP
GgnRxDi5T+Nl6d7CziOoA+XXPZhtAoaKhJnHmrC8R7GDHwCGsoP6Gp9FYs9+hvSF
mE1VKrVkzpjSa/hrR4dmqS+NlRcdlLn0OOxcphw3UHOAOlrEj/IwacoigBMjPLwV
Mfo5DjHgTgK1QJ99hnGefDwLAXZVdByv8UMO+R1TGcMz52UpQ8rVjhYMB1+/Q13e
Kf3CWXhNb0vGIcDd5puk3zAlAZorZ4ltwtwO095BJIPPmw7tbxlH0OftUNkmDN0F
4NnufimuDHSxbVv3ZXjUW/4bCmmIe7g0uJgUdutQ0P38+3m5RJvdY6YFcttV/avR
6p1ELhLD45ljzKv6rGRq9RTzsGOFw+vSb0CRm+sl3uihiqqbp0Ew6AZYVnOXqoD3
ZurFNZQFN/h/hwj/D+Lf6yfa//reSRVlemzn9xJo+MxPpzbrraY0EgKMGzopS4T3
cVc963NnyBboGSz0jVGVBfie4SSxUgTE3vNmE+M7r+/mg5OYzjNsIyjLPz/9DeYZ
KbgbaDx8/Yq9ywkBuiHG8DNSeJwHgAWwhVxIWz79bfjNsPT/AXkTkW7hOZTIQwH8
hgSkrCQ/aNEv380kGZJg7a0bFWg/52h3+Vy6FfkkZ2zXrSsso+FY28I7jDTeT9de
TvnWivJFGc7FGCLiB+2l/rbX6BQXf7cf1yzaHchf23WK79nRvkgEXrA9t33Z6Ewa
oAtCPeDTcJCHzztu6lSKWYTiMu+Q0h2Syf3tO15pzvrDVsqSkVVDUm+LRM+QDSs/
ni70fLdH8DmcWoDZHnmKXHuJj9qcAGLlMtA7hW4683a+VYQVJfNkBWc2lvC59IW2
EnwV7+baXpOzkvuD7pPU9qy/ZGpLK9YtfH88Px5rJuM5M62/elYUdQirLm05Odg0
h9ijEUsygqTPczyoSDgpo+4Zo1b5zo1ElC6Qz+L8Rst//nQ59BS1yilhwMJBpyk4
XkCQtiECi8YIU3Dn3v6SAD42xnnGxQYelUx3OC4RcyX1FDxCWHl+8Qs6rD7RELp6
phGa0YmNo4uNJa3to+ddvYr3Q3oN70ckFvmbDm4ecCW0kWrDUV5z5UAKU1RiUTHz
HIe8D7Df81B6cV3cERPCd7uA1txf3ZLaOQjfdZYJacOxl65xOSIyFnpo/i4xWBBT
k1nw56N73ACHwgfOStlyYLygL9pGe8hxYr5tVL3kCyQoYAg3mVBPy9h6qa5UCA5O
iwT1S8h2JzjtEyDVAIWEKYtVjGCY1lXSJDfpjGieVuZqDkO8YohrUlK/zJNEjS6G
SQPraQ6oxU81pIyg8u/W0EiyMfRveUll6DM4DO5Jl7xNdg9YKTIJOgX8p2oLpTAI
+KffSZDLcwliKygsl9fsaHxVyVtFWvCMUnTaUgvdS8gRW/Ns/DR8pih4QWO5vO8A
3lX9L3lCBSH9frdFwJ83M7BEBvVvbm0PsgfAptlIXkY0xFCQuf+uZMsJqwuEmhCo
zEKzDMaA1P2OhLLYPvHa+Dd9Q8vKlD4W7vg0DQbNlPNx2UpNI2rsx2rWHW3qGVpu
3rZ1UGz/dKPyop3QbOtpylEGALJYkQpkeVkq6WZ9gN7cl33ZpL7hjTEYoalqXy+S
gW0+kLEFX72OZdLOwu9NrW3jG9EZedoY/fYCDF6nV4JEu1scFaFebAtjNtcQw32w
M/gXhQZKMDZlwce7sc7JKM3tQbM8cCQS2P9yFfldjzXjoxwtPqo/YzVHhEL+kd6A
tkWdz8mtxGHX2AzguRPPwPlA+ShFLj3Dv9V4MzIpCUYfJKp9NSBNt/JMWCFShXgs
wRT7VgsSbFpldHjAMvGwQwon469lGxq/BpDzXSbz9z1zO987Rc68sZwdc7L1wgPt
tBqI1fsP2jn4c4JmfUyX8sOdxiYYqdm59t1nrttHgzKq1UK/naWifE84WW8LUTCv
XySwt4Imx9ZeEWPG5QyPaTHEROp9n7WRkMHK9XKxUGMdsLu60MU/nyWOGSndwgKW
E34p4yzk+MhlOYldjCszQeGmBuv30bizrLWbt46h6pTVuyjxHS57kXmkaAw/bOdb
w6DkM+Qap1GkEVZ0nnpijIsp8y6abrYoptT1kMUxdv5asrryUmtSfPuYddOvr3pg
inNfpdigUm4uszTrs00E/cpb/6p8wDUDSLIJY+YXfL+EKgq2yB2a5mVyEQAq68Kl
KPQjp6hWWmvRtyECDMckb44vPdj5riBrc7uRTNRAPXKHYnQfL6a5flUMgs0cLMy5
184xbh0kPTFFkNfvK1zrFMuMiHpPvp1shmw7CaGoLwmLrPnv2K4vHx02iJRUhtlW
ouPFNoQO7VeXl/fOl41mMU0iXIXKAlEiQeC2agjyt+jCkA0SlOuoea6nawSn+Vni
nrBH6jXv1XGipoiu0nB2YxSVF+XVWlAClUj2oDMl5ihs2qIwq1Kiit2Mv9iBWsqx
KI/nmoZO9AlfBd95qiC7GeR4PBEzRLZjCkLOY3eUxNF1x4VGK0LndmmhxyaYmg2K
v8LlRy2p2jTdEdNnoB9LTh3LHKaMkvZfDYmt27id58rSNeWC2l5Uft1JaqzcUe7E
6/xsRJhGDwPt6PfNuxUX2WkZeIvauU1oHTAxjt4BVsCRU/I4h6H7AXdpU4K7VdDR
HgON8uW0MivAUmt7WHlWSQvOPrg0Ke59cvFRt/UxdVzWgz0LWQp8FT8KlXrhNIGY
Nb3MPnMnmzIqPTNFuEVzcJocKuLcDsUVsZVIv+k6t/1RsHK33tBZW/3Pa6mrs7nQ
QIbyWV0sZZp7M+UsGYqK5byTEuWULj8ikUVD7z943Ubx3dREn1TW+067YAudK7Qy
dUavM0lJvhW8AgoWz094abrmWndQ+8GhgeIZzDldIE+TTnqUh87I35rs62fXdb5A
6kIaeOAeh1CyX2pmOKWwCMf8OsYerw7Hd/zxpZvBiLJKmYEP5C5lwQECWHQL3gFZ
xkY7QjamFwXpWLkLIOI3sZbI5GeBtnr504vPLQ93gyf5XngYHHIorfqmkghzaGfY
cxDJFa0/ndCkiHKJVliO2X9yLzYdwzwBKSHgG/JcXRk5sbMsTs4LFYpflSBbEJ+8
bFdyu37ACcP5/Uj73x9Yfgl5gsZ3lZx9QtnjFTqP7xmyRvs1xfdMQuv+uKr6X0Sk
yCQsDrWmw56+CK/YBN74GYKy+cVWMA0LYFAc7ZTwPZIId4J8aioDoy/4u+eCwNMp
6iSDmjo/4vQ0BkLzyR0zo71oEZLgOHgmIvn1o0IdPolNbI0QElqI2ChjqFz9ecsd
UA9KUrjHMLlLAFlYcMZZMEoNMhH7W4aBC/ZS/zBeLIFEL5M95ZgLq3tBGLdUyCcY
SQdu0WitT7VePFswk/a9lhTka1xPwePJFC5yqZglCWedmTjBhFls5q96QTti2QTg
3E2vQHSXlNFHmPn/oQWPjoWLa8VVfCGbnLHxjGgeXk5evZneXfAoZFVxRGFv8BN4
+PIp54dZK2WJqBy6wIwlngamB9HImF03G8jdFBJ/rY4FRZjHiM9ipyVqB0bHdNPu
CxkTQxXFVkh0wIAeNm0ubt9wXh/U/1G70jTzdBjACnyRCwATt0mNDnvh16ViDIKZ
O/cYT3jfJDeUzmN6RxpK+58/IyOIYGwl9FrWEm9+ufi+QhhcDxbTBmOI6IZxQZ1V
Zr0e73gDE8kxliTOkyjQQ5Ic2kcn8N0wCpIJjMtIT3wGBPwHqjXkvNGJp7asaIQ8
mTDkRmZWgKN6obbvnCi4Ja6M3C3BVXHDcuFM5RVBt3hMQwOweFt0tBeIOaMW4xO3
8bJ2ajaVO+9g5idJ6nagbYzBv/P211JnK5cnBxQlO/Ljms7S6ittdTHQRi6a7Tl9
atnUnGBC7++a3q0TjRcXhDC7Gkfxy3fUD7A/VOUONQwhanENWvephxBCdUGw1mEU
/xkxrSXiEcBBjoEFh2qLuAfLQUVJYSxRbMcJdRLv8yCGwZOOR6Um3Jx5uFrIrYFM
xj1BhxmFEiX8EZmZx0OGaLFJq+ZcLE00J2lR35nTCjXfqaEzb3nB7Xdb1naEItwm
bTdEWXQ1pXGQG2N2L+JpqJcbUIYl0gLK4YiWI3jnp4SJEbCGX0RBi288/p0YVhtQ
GJvAs3WN3tKkHxaZt7GkKbyjvSnaqHFO0dEtaqeboiwx9UQRDY/oYAv6x2Qm3il+
nizv8rAjgihzt9CAYUenxtEOCRCicFdoxtduC6Rpal4ueNtkT6M8GDjdY73Kza8+
CwE7/5wMoFMYkrHMaeJzjUR7kWQ4Kvks/uOu0y0HTYoTQ2nOWd9TIJsvFtYbkXXG
9cfrPRmPoqCgCE4/ZRUX56PPnzJ4YiOkziJQC3WgleZFFjwZ3qqp+LC1Uejn4R9h
HEMDqU5Fs8aQ+rLhw6xViSzN4lJ0f9J209//XbzdIP0ggd9Fxom/DylAUcY/M0mO
Rd5RSkmC/EZbtS//iwwfEQBqG0Pb7q6LeKZuTJsvB+Nn1v87/XMYATBhatKU0q2C
eP/e7jywzbpf7P5XNxJoxIDWoZY5GIO57QGOH+cJK8gYWcVgPKEgd1y5h3fC05qf
C9k86tpCTnTgFcfstr+kwrG6sM+XS7ZrDlFx8HdkbRHLc/nYbcLJBfUF4OdTxA+5
fvSXh4ymUMq3xkTtte/NShiirszZPm5bke4vjmro9ETJDgj31Djv7pneyyvHzwPl
QpVxJjgMpDQVQ71iIy/jc7PvF8PRaQ+b8uBH+khayJjAZ9ZNslhky7nEbj6mtonS
Okt7EpZllSSofyFv2yJC0yCFk6bc8LZU4oOL0yfaPmNCl9ZoaKCWclWaGtGKmYtC
XQzdMiwvfzbKuwGTmEhDSw0lH6h86UC5QhotqJhLsgbak6GD8SilqGLj0OnjUOAt
Y3g3qCMs2fDKOZTYGaZRABHpTQDv8+Pd5oMCEnc88KFa9XTzhn20Plr/pa+S6bnl
Y/xk8KHNdXyaEZdUUIxQxpO2k58aLxbnmRalAh7adXk1PXhCMSKh0HjabA3aW6xz
IhnOlKH/ZqUZ3A8y1qBWtA0P6K+MFlL2vuOPl4rhh/p9JAbFH1oN5o25CkuZB8WM
DH1Ev9rzsDkghawZMch2Srw7LcVkF5uaIcRtfahQi31EmGKYJDlM1Jzt8i0DO4ek
59f+zTTW81IMccHM8yNktxmHUwp9saFe1uK8LiS6zj2B2F8tx7U7AEVFoL81azOQ
ht70xtTvYJ3acM1+B/1T4r8b+Vem1jvQNSKS9YZ8JjWBBgHjxsma7QG6u0Th1R3C
OCZsIXl82FfomSiFqABGDieV1wZI15uiE+Hy272+jExfx1JYbcmB2Faqc1GDnra/
g+U7GU0RVMamvqOcdAMB4ONr8KshTCaV2+OPEyuKUR7zHTeLLxFt2edoFk9fxhW3
NgW4LqVWnuShHvFrSA91+c/+OmfSfdYBbgYOZVQbGgg8P6GMM/8qtWCXNRLR1wSg
RSn7j3JnHTEVqBypxDq6yTLWrsmoZ/42Gxrw5Njb76b1Bk3FRTb76s7uBoWjXhpf
YGhgbLn4YKYLSu+VUvGq/zLsC5unhpMHgVFYHHvEIJgwO2phQWN8eXsgSifiBI53
uHGn+EVwJpXwcKe3dAz9QoRv3l+JlS5rYeHjwnvQkJTJrSSlA2PiC1eg415EuXHo
ZdKu2nsxO0Sle7kokFsb0/3mjoG0Lu9fil+GUEkbXGvxwINrw/47EHmfYfA/VEP8
VBPZnLI5xeR6idjL19H+kJPwVZZ5M5i7BnVW/qvu9E6uJHOX2WGpaE+FaxdYhuu4
7lxV8I5l2NguknubMRGgfZ7FhfSKXGS1GXnFvd5xu8pRARVIqJKzMkO3aamE0mF1
8wgrQqzLaLE5tJxc8YRVGxVYegEHKoHSEEZQCJyC9Erb/Hxn74owAd/LvOdXkwo2
yR+oWkIcwZnyaFLGD4fPecqpqqTK+UA1HJx8CzGuXa5FBNxLOq2qQgkKmDuhBHXE
od1wdvfz2iQSyBxt5gNXgkDGM2Mff5FYySWIHVlHaaPOkEF3SgTMt/Ipm4E9yxZz
yI6GXgjyBq6QJa6ZBvM5hKkbtUKBjvoR4YdsxezoBRMFlBFzKwNsTQgenOAhmmpY
JWtBBTzJzgpcQVjZnM2Kdy5GLBrCP/IWjEskmsX9Bgy6/RwT1x0EbtFI+dVpkrRS
vdGW6V5+sY3LALAbSJ7Yj3GLCX4B4CKoKTJ4PSk1fLF8AuMZWhF8tj2ahuyomWhm
VjQWLmIzqcIbkYBNJO9xM5p0wEjWDhQaSb89p9aw/q+XpEWF0mtvuCOWkfyCJ0Yx
spB0yYxsHh7Ds6XOABBVlg1AzFN5d+5O6f8JRO+XHdXlaPEVT/HWE4MacR0KOCnv
i7Zbv6dMfZy5RigUgLEEydrFL9UShu6coqXc8+CV5HSqh0qkcEs425XmEgCDkmab
49LlMnwbKlmn4Ngslz5PEOoRmKmKM8ftBpz/wpGtb+2dFU+keTs/CO/bvn02Vjee
X8BVj7O/CcnrOPdug5PTU/HYAB5r8WBawk7tNfzHOuat7vj9Sa95h6OqQRQVNKvd
uU3x+Rx2OHhnJr5v6Z1dto154n96VbpEpp3W1uhV717J7YNIYuuPyr5LI7j0vAyr
hgw14NDYJHxwjs8JeCH8S+p3zn/oYoJv+StPhduyjxxlClNp81xuhKTkyhvEDKkw
p6RIkT8tZppmjoKxz+yzOcPq/wlZ/AXsv/Y2G1d130X+3LkL1KskM/xnAU9Z0rwF
+PfqIm61DCWOJqMa7tnW1lxXuvzEQC2htB6K5XOlfJbkM4r8ZL2ghv1lUU3o+ULz
8hWx0qBZLCb7i9xgWlWXPAq/u3LD7DGzDKJhEi8bGbKn+tGq7/By2Qi77Sx9+JIA
Nd1XjQBXhfgAIxn2twHQi1m1NM9S2DnOkyu/1pqKqQcTk0K/tIKDFzbVymaWddUX
kmKhAj2HDvGkCXXmdqELgwKZW+fZLN9NvZLVGuRxF8cIJj1OVFPCRhixmgh2/nim
NDOiUmDj+o6R4VoRq0Ytr8W8i3i2S0yN4c/HnK4bChx2xHmfgOI2euXkWNd2IqRE
THIzK3ZYA8wRcwixtRnCQpyOH5fjy5oiExiUPqdjVlV2BtBCPUm6CvgyGFHdyvYK
KNrMdHq7gm00HVhUXhhagftEdcTJut3p88d0XML7slPNx0O8+/5adnD+cKwbt6Bs
sG7BCtYtcNKyFS4qVl55zU6W8rnmkqL7EhhED5xvbGBIZ1fmUusNb4a5ppC/Q5gO
id8taQJx38/BDC03KziTpHKzFaR/RHuaWj5ndSPPJ/5BEd/4E4+OCJGOBkMY/wcw
VmGbddDK6PkuC83oNJoNNPjNIkikSTdv/DlpAeoWTTXYQpPTIXkQn1P2tQDoZZnQ
k5DcGJhkN8mmCw0CaEZasA79QMmZVL0uvq6yRqYh3jEOB2PL3BAkaDZDL9Lnck9L
4V0OCLxeVV5fWG1lc07flbuGLPXashK8F7dQ2q3WZTXXS/QZ4pSiG0/9UX5AoUoe
PDgFJsoeIAnfYRQIK8v8lmf9nm0vXlxq/e3JubXNsh6M3TRUh4b7F2yLlNRUYMZP
msuqCXRyITA2ZKo52/fbucwGu6ErvLTWb2UiJ4w+bCsYKZc6+qLW2os+dFzE6nl+
q4pjUqejimXu8y4QQXOIgZHa6m5yhqsSPOvaqHJpQf3ro5OX/piGlMUGeMwJ0SNl
QAU98ZUWxjf6he2qsU4BBQTQBBNBA/P1hhm+xg+De+/SxWuiMcAer/bCbQDuT0i7
nUsFNG7AkQPys7JvEma0VliumKD2gbNkfwJffOuX4+jRqzSXyRu0Hy/pBUWbmebD
pMK0HphoQ/icXlB7qirI+c/hikIzr9bAbEin5eHq+2aLeF7QDskAruDg3bkuEioM
yInsFIzBGJe/l80vMlfJaU9ZR88qDMSolif0eI7thpmLLPhMgmyhUaaRmyfTzCal
s4OuB6Q7eELz3BnRsGM6yr3xqBx4ALMV5SmemUOJRD6xUF1vlFf5RcMwcHhrMoHi
3ek8ze8cHBR307LAxhrXiW0+mySZzY6JsHanM5bx+TEJUrhMfHePzh483Jdguond
15rnmnAc5AWj3sli8FwMD2rqU7KbOMgvucYP+QVNJJ7BqfB0KYzQfu2FpjLTNO4u
AWjScC/mVsprqoSmc5uGtPH1EmTfRRnZlAg0U9aJ6urpT2HxWdCnd28XivqhB0e+
w/HHuKXzsjYSmnLAI7hwhZgXiG1BG9vAILs8Nqu1HA2Ex56hvVoUXigSQthatYkH
WkVN7/pZeihlV7RdWvJFRHlo6O6fagz8wQeNoRHZn9OyhJJ+L4Y85AYH3+2hfR3K
nX5VbjEPX8CFzYiBWT41wsYBWM4T5bwCkfirMdbAKBFtx4rJikQGCG5evgADL478
Jw5S+M4yLR8Etixqv8gjqlGWZt8gnsx5qEqjCptLKK5MDnGkXkkd6HP3hlNLAN37
ERuigxiAZny30b8Ahe6qx0dO7L3S9g46lwamSKJC1BxSiVsq3jyUTkczNaqtKkWa
9+d52fXlQDjgZQ/kUZqarU5p6HMjNkLkriPzMz8EZgrQkK+mKFy4E8DYdcOHV4C5
6eDzC9W4UmJSG75AIjEGePm4NP/Hj+eygrlP5wtouFVknGYgrq+irOpf85G1AIIw
Ht9e1iAGPpS3v5iiFl52iM+Krpz/Hhz1ZKyWstLijsnHf8nyZIW+jUgrx5LaADqF
tPpVcwomquQbMtykhPEG4hjaQCHKzIS9G/FHP+rFiVMC3Sp0EwYlt2npdYyGdxqi
+K3LIA/RVY1I/gXChYbdUQ6yaKHJJJ3c5nAy6turHdNORlLUX+EN/Vq8Tg+PsOlX
hpK7+2DgyWKogdi35JcqtebZ65E38JNavZmZU/hN35vY3nXL4wqVYMjg1B2m/kmc
NgspnpCR8v6iHmVmSEL6stYwX7iVprsCSrr46ORrYGsOSFPLWuyghxfrN0WUE8FI
+EkY2d3+95zizw4ixEIsorlGNQCHO4u89BVvfwrgRkaxkd8i952N+GVMtCiCUM25
6SQbkmvDzM4oiu6luT8Iogu6chUGftPtKG591aVHbFYDORUDfyJdOR7XOxMnuSC5
zKo04eDAv7Ua/+x/q8OF7C1u9IrMUEWFTtAHMaP9DDST4r28GCG/9kfDaYdrp4Mi
hNAmLTjr3CNhpzCmhvM9NfKHYpnPgNGO+NPcSAIH6T1FL0o7E4IYvpaPtGqerR6M
QTOIilxoPrege9fVYaBUS1FickyQxfE39Ifpxth0wyewpENQqt+8cNCaRsGk72Ji
ydmHznI3yaOwxHNrnFSt1LQ1n7c+e0cHmiwDITucZfGgJwILZC1SOInbVPdqzMym
U2nQYm1UJ1/VelZMtfL8zou/YqzuR6h00YvSwxMWBbvUpBzOguT01QqEf+82Ic07
si5A95UWPylDxwsFhgqcf1G06MuQZLI35shSycCHanU9xPLfnNkL+2EMq7C++A7E
BY2TMjExHJGem/A6H4tNPRTp7pWyKxkHykDvqHtPUYGmTzS84+xtkK2ppIz3Veyi
7dzUFyNPH95/Rmm1By18DaXMEcd34QDCjtt5KGqwEO6lZyiw10yvBz4V0jYDu4o9
e5Cz8Y7g/gCWvExWBXTiVDn3WLAfzo5/LVxzqM7XeMAYbglqQVlLMjEdLIccyHy7
XFXmRtxc7x7Z7ou/uiC+tWRMhmI3RWqOqwJkZlH/MrHCE+akYb/ykFva58Pntgs7
aR5K58d1gLAmg3xnoMWtbMIrk9mXnYdaP7w34j4uE0Cw7XSkSdHUo2tTp7CEDJGL
6F9aNsYYdDtXdF0XR6PChIoeUyLgswJg15fMBEYK4yE0nCfXiPML6wCxi6UfY3i9
dJOxNya2RV7dIPVFJMbYuSfr1HevfJWD5uBYi0qV1O8Nv92yLMvPWnN4ldd2ijs+
o/Q/Kt43ZjKaOr40/zm5byrhbpZRZm4DBhjwtQ9HNnEykInriZYW8yyiAINTP0WM
KJFaE3gwDjqdou2m5RMhZu2cYigT0/uIN7Ch3c4vtcTHupCvS8pbnwyjOdUbyh8h
MP/BF8otylFRILypXDrs6jv4LlxDHF2i+6eSJ4UgrtVNTjjrupPPihvWo3Vsb2eL
ar7yLpH8yGCyTgBLRVwCvt6odsY2NjTMcDpnaRZIY8k9kIHJCodIU5APCbVE772D
FBsKIgxYZeTKz62vtEIe9ITAXf5URfBgf9EGbn/jtRCumqcwPzK4MqnLDmtvGHHe
lKHhqqIYtvrb630a5rERPIIFTzaMWQtDcLiNxVrE3i274k/ieQECn1GNB0z916UJ
pcikCHzcrfjl/t4YgYaztQZsN58yaO3oJfJKnQDXLLPPL3FFC3qmQW4hpX9Lut/3
YK8szkAleDHlDgi4mkM7J5yh8of3vzvtPK6qym6djGfMSFm53lYjXnibN2kKbPbN
8bIRnNq38dTOHAKG8NNdszvWsKx6QysaOeqYUoRaQsToV+5qb+mJcF9C6rmwN57g
z/0oLDZjq7H6VZhjPIcgnG881GL9Xn8bPRSKSjqoqkpbpncbXzRj+hbLXOR1ZxMp
lfM07Gqk2ubRDYw2B0jJnXax7uqLENxe/CymKjHLt86DZ+7I7XqqPnNvhKbAfQ4h
Pwu9x9/11XFEc7HpBDo58YJKYQvGkm1Z1oUWxwF0GkDkCegbr2dOOEx6eq6pFDee
6wD7jW51glzr3QCo9a9LsTpQXNq0+CojsD2dRy7nHxCw97RfPmPNXnnrl+TrLAb+
H+Ryh3Th/7CRUvUf2+ZdClx3wPkdGov2j0efbrxiy8k8fippcBW1G/pqWRkZgkz7
+BnbYL4pAHAGJ78EsFCPoSDTnAJVaOsgzMrWLDUT/+s1FV6P0vDUCopn1dO7g4XY
XZlk8e80avSOxv65virH8q3VJki5fGa0vdiV7Mwwl3RIneGvbFlNn0Y7Sh4Hh/Ak
8HADgvkYiO45uipZHEQGLEWh2HeNKRhQaI0cCvRmj/ONkxOJHDycudIuou7ZjCvs
Evhnxkqhguu/SUXDNQWberDSfdphSdONnZhsBnx/p1uRS888iL/EYE2NtxkC6QHd
Z7Sv2ipER4bUeF8XULWc+HlwhEZSh7iPAPRrxHJR3c/4ypUM/drE472PGHFo+QU0
Z2wb4fJ+nbvVckF+/nnASJz4HK/4I+rOyhyhNjRm1v/YI4P/d5JzFtxoRnHHrLVm
0++XXy6PtjcRcJ+zTJNCxMBzvzNhwsxTtl4PJIwPvdq7Qn2siDIByj8VDNQkKNix
edZxXcCmBOj15wLsolUeNs1CtUIK2Cv9jIG/zxKDfcQAEaNgoOcGAT82YH0vpdY9
0GQR7xp4JHnIPyBEA0b5Ox5f9JVu6i+a8PQLBTL5Lwq4uEph751P8XB53QMz1F/3
cVBl9eDa/vvnzqUE+sQtN9jSW93Dxo6P5XW2txd0VzKjnoPzvRtwR/uBWbCNfJs/
So0G6PWAPeJre+kOAhQlMwpht/pdVIwQDd4OJcWF3EDHcbd8/i1eiWb+seTteG9c
wVXQ8Bb9qomRf8FgQLHKh3JXw5PzPySiDOONTRJAuyd74n9ZvWW5blPV2uIUYkwV
ONPh8b19U1/wJ9rMOuc5IKE1sILYeo2kQvaL1/HWat6vQakHXK31g3bvVG7L9Z0W
ifa3vitHj7wR9M5yL26bXhp/nJKNjrySXizqeJEkmb7qOSsrnBT4yzSxlgQQiY/0
qo5m9J/R0VKRraNxeMMDHWViKqJcRDgSiY7G292GasCXShPZvuVAJOoZYgFCM40w
JkXnDOqFMfh5oJlEG4UJf2Xr3O44Tm2TqZEbnr9g5XEaYsTOvtfTn63W0Z9a71jU
g5MjLqesEb9yW80Q7+rpSQaHOQWAL+Ie25IgSW0NG152KYKUycr7w0D/+c1lseMO
s8XFndVk6C7ZhEkyecLrho/ZedcTf8xVLE7N/ARYokbNlT6zJEYRKDMhffb2TR3W
a0jWUhCU03BvaXA6tjP2nsfLKEv+KoWHBbtj1VP0tUFNCnXAtCq3h0Y0nulOCuPx
jtDjnmpWRM5SMesb//doNFxFM5vTM+TJ9y/YFlry96dW2gm5cPRA+ugDmxBGoRbs
up+JYlvMacbHC91JfIftvIihEokWVbSJ2aGXd0UCqrp1t34fBW//P+zZjlt6MFUf
VQivzQ9/5GYbINqu/mEt4HO/oKdUvIZ9vXUjr4pSsliR8ny+xYlNEOffXtsEBswN
4KAfHYCK4Sx4NvsrzsEm/IcWLNhYaj/JXt5ixWdtxQM7Ygj3i1VDN4ydfP/oxVnq
Q6P0gdQQgLuNJZXCwqOHq9xFLf0REzkquDuvsTuaeNuJH0tQSPBqaFo4lWZCkegR
zCHiMCqiS44CziGglkDl3Xl37P5OBo9g8z5y3Bx/UkPyu747DgxUVmmu0KHuiash
yCOE5mI1LnqnVRr0uZwIWQZrZB1f+jS07HXaJ42jvxjB68/IRh5swxraTjiacrKu
uS4Hel1zcGHvsDzljQquQpFXLAo03UgJQ5KebhZjaNdf/OrF5K2UJwbBQJPrH+RS
duuXRe5+g+nDfRn7D8kk7ZVXj6HpW4PHrryewIGef7NtYjazL66eqStk9izJniKN
c07H2CAZqXcIZ0f2EBVAe5XSENh2oI+HdGXNrQmXBqyPqyrOXGprW15keMGPmVWd
pKu4uU/A6fnZdQjwCEjD1E4VZyAVtmrOLibrXimTBFzQ4m1xstnnJb5FqU1npvZ/
BIojePvVU2/yJGfNuwad2tv3P3vJ5jeK6xTy+7l0LRhGnd0CTsHjPj7WogzkGRRC
tStZ+r9KpJmbzTfXjPgmjC1RF0a1uwVhc6V/jCt6NRenEEmlgrq8XVTCCbYovqGp
SKNMcQ/SO8bbbmrdixbitFRpXTqOMcOZ4XrjnuGZt2Ju2clbWy7/fNvn9awQdt9r
tTB0ofQxJLq5Keq67q31PumxWqjl3KDWhonGi4ijRJJ1qSDlH8C5shbAnB5Yn2l7
mcM0vMDUmaYLUC3+o3llOykzIrBaIbKvJYxiYyYeKcTsTm9YXEdpYQnKPw/9s05R
ZODU17VVdNtuK3M3SbHpSi8VczkC7tIhw0Auftc7Yvum/8mDYJGANVnIzM+hV81j
yexY5uKtemfgn0k9u2ndI7aAUMxlHJxuGYJN8CyOl+Q8NKrP3HyLErapOGEk6C2s
qhNJJ3T2tzCeckki0SzH8Ehr3bLQH5inFTL/Wbr+NDuuKe/TqLX6ZYqvvpXaiRUA
UPx/ABOqy3xCmH7l7MhjQYiL36oLdRuMK8wiVDZCkPaNJ0j2cKSHnXsLGANugkE3
Eq7Sdn+MzbZxrhNaAD/cyoY/V4ZbOLu1vRzJbEqegiljr4yA5NCIHDeMVTgwjUaa
0dDGlxt8aAHhz6hxlXza/zdk54Lr2o3vutB6F59z9Q+rci0AYIIcMq2z7Om0rwtd
dNknW/5uUacR9sEYWVMyDUEfd4Yed5h0tGbPYV6atlJIp00pIz+XzXsg4QbHeZFp
IkxTneFuiVuf5121ep61ltCMQ+uztjWkVVIBjZjPFHhcenUxs5cyQSrfbOTpzzuZ
iFPWxNFNQyQcMK5Zol14REdw9QQUCg7+DfURcQo4GMhQ4tmHp+A+qM6eEUcw1vEX
YzRhvryhuRmaHOFaVZxEavbGDoGpaI46sXSirBcaJEKi90gnqsySSX+Y5MeoALaJ
hlPNNgKswuN0YsMIhCkOVI3HUQRAvW+dZcK4KhsCvTqTm2BtFRLbXMQCXIg+85LJ
xj6Mrkrvp8tUBl/80Jm8mSHSY3qCdiCEYcwq9vUNn0tWD74DmR+Bz7YyjbWEz//4
3kN1M7bXl3yives8x8j3ZsAKh9KVlC5jTmuiZBRar84r39g7a56Mn9dBDg+m7DNg
vwEfZSBh20O1geicY3ybWQ4sxo+4mB7cf9PC977grwj0EAl0Hz6qoVcRbnwE0rk8
JUBUI3g4jfkmD4ohIeiWXYDwEwIk4YIhT/go1nfHGT8/5Sor5pYfcTJ2Eg4KX4th
STAPPR8iDn0VsF3kOgreUhIwEkV3rh627hN3pgkUFBM6Lqayf3LPNfKDN7D5Xg/x
2y6+aPtUSCjnEkgKSw+cmOkYrAKi/mkTksw+YXD/wgYz5GAVe+XUhPjKA/ok8Gxe
4UNCjfEq82m0PnMGpHfp1LsQapRAedCQoZokOtQKCl7qXY/TuRKJcnogqt2J/Wba
mv3tnthqBKCG/ydmf4xeMfSr3yFtwCwunn61K8d9dz+KxWMHLSajJGrYGYo+CKA4
JdMja506EmMd+7L53bJ5/EOJDyh2TAgw7sB+3Ny/sDwzV8Ff2cYcnUNFh3hw14P/
1ntvG32VCdx4Hi5vj0Dd05xE6qe8JOT5fZ+9jKsOTE4FbQMVujcTYB8JUQRvr41u
yLOOdw62WO+SNl5m4bmOXltKyvPKkju+Xtawr5OuMsIYN4ecQ/ZdfQAwdd4790PA
gXcNOiB5NDeQpdlAH9fK7LACuAyaeicIDVXhuO8oDPKwtKV+TaGrOQV/4hqt4yPU
rCTrJ274msFpHIMWSFVXSPoQd1oRp/EXXqXz+M2QQwZPg9ZcfmNhUR7ymuJtjbQS
HTAyr816qt2uLbeafmL3wGQhjDqHm3yOgwUZpf3qRmJIZLm/XF/7eGxXiYizW06T
mHZ6JBwxPu1m90ga0XMtilNP4b2devNw/fBM+jYMbHzVSWtJ2ABAK2euAnEc/GTt
srcRjOAAIYQsYO0FMFvtUplEuJAPRUNjsQFPPMrxWoge17yih+ADmvSU4HMUYF45
jS8b+XZ+DxPOR3Dsqe5PjkJC3JibOl5wG25uzdXHIpA5fDV/cvhogLhgiQgcwPkT
6Vy3Ob+6easMMJEsS1xXcQ3Vf0sxwKaqJ7Wq1hZvSJ0yyhGFS86VSgPmN3xq8WZC
TXH1e36/0ayYtoTUpJBdVOELD3dnaxZGBTZak6A+zSDAEmMu3Rivyskt5M9WChv2
iTpi72fdVnh2anA6Wn7DPvn9R5CV4wb5nUkKHcI54AEsvkEmXn5L+6z/Iq5SdCe0
CihsZoDyROdhk60a9HgVoW9fmTg/T7vc3DJGP7cMi20qtetR5l+WArAWi8fHVBfG
zqjDNA38uW5wlmQTRqA/XgnExoH1udMIej9j6pw1o3GeNkjdJRzv7O21X3OODvd4
3bFA18UqkmrXXUVLMwe3w3F+TOsnNXrrTvrhQVZOt4PNuLCHp4Gge0DFA0xEq/WI
WLyovtd7wtwc/QJADaD6f5o67SZu5iRhuwryQzeataS0Fi8KBW1BVhIqh55aR9gb
PhrWg0i1bub70WxrbnG4pISK/S3I0EWsSsGXMHbGalLsWj0H4aXQ8pX+Y3mJb7At
X/cAi+5JjLBBZp7Xsmzf2BOvAVxFizz6A5xTd1v7GK9ZQzs68mbnGMXRFtmDECL8
aBQsPGYkkieIq4esmTIwavWjYbCUnufSTGRkqy4QpeDx8QYnfXyhR/FBEkN4sE4P
ojx3+1/sQeBxbR0Tw/8LUOIxaiZT9tZB+1UQ+QjXENf7MNcXjU6u6C6P5DehJqok
o87JBoAwLXkVUNrYCupVV+/6y/sDSX0uzQO+cha/pUkpS3js+mG8+eUpZ0I6Ty6w
B30aGS/8kiEcpearVVUQ3OuNT1Ujr0K817drkdQ2zJlvuQZ7pGpVO1ewxJfYybGv
zVUUQBwxgKkShNmfgaHk7sUJccGQ9TiM6IlKI9QvpQd3OQwg32D/cjWX7BvbJNse
vyBBjooaJMiWtyatTyyp64uuvZCePyQrAtkUnEn7s+7AgyZgPBCFRD5/yDtSS/3/
ciVcZkw0XVqstPU4wBNbsf53cKeMVCxGuMOCasHXiBIahWeBVKAiDGBZrAdkBJGE
hNdZUGP53MhWEjd38IH+ndQcjkPp8FkSeOS59N2zxhKWI5pWthaTAs0+9QLfUVvD
xJgi/DZhr6Qqlm5e1xfx6gFuNuYpyw976C/13Cy/kGEWRbGhtopvbzsILr5hHWpL
KJAx5RFCpwZ59X9/fBRcCias7xlviEWqZxdj7Yt4FnOIaORf5zcWUAhlMYeMkZSR
/x83BIKzh6TprQGPpDJKPPsX61bsnZoa2Vtz11afAIhFPYLLelgtDoOizGbD1eTo
Bq1MENKaa/2ze03JRnnWLA2IX7E+Vg4KEjRyeQURNy+c5QbvcmiLGCLNghVYEEJJ
2HbIKyKZw1YXXY85mXC2mhkDD2Ylm11YADN1FWnjMCPAdYZ1sa6lDjoVi4rU3Cnp
w/y36GQN52xXZgJjr8EClowB9H+hEXDXAaXRjrerHvodqc6vLTFCbeULn+kdONWj
Z2XNHOUHR3M5iBTZeMcnFa+MdgAqbh9Xwj+OTKyMoTSj6m8rde31ZsFFlr+aMHNa
WUhJLfbyKTawkezVWj+YI7HTQQU3AznEMtiqAp0a+wjgujFoNlkxRpAydwplUhZh
QhWFG8un5O5vcHWncqbEcqo2pVIQqCq20H6DeNvvxhmjni+HY57mLxCWrG+vfxlK
o0xqqCQeDJM5p0YseX3/orkeEs9UCrPefn3GIoDZ0oT/lmgnzLjP6zMmL2fdqexz
ZhRWGvwgAcVf6PAV1kC9qfCjz18pVzUnn8u1xMmV3gCgoEnHXIdmp0sdp4HUI9Cj
ymbekTHOjFWYK+YldHnkahEU01mrolo/WfTYdGB68pKHG4IrCJc/hUS8ykS5fvT5
7LCsMeBgbP+RfwODoZlSmByulahaJ9M6WuiaBkSOY+P93VvAiO85zaWBJ6XbJlwO
Y4aGzgypLx+ByCbLJHuGPF44ZfmSuMB8+P1tfUiPlIq+vYNmWbvxB8Cw+VdkDvEb
7/J5p8RZnZZjqESfNasRdbwuBw7Mi2eAHVMltAvFzfrpSabQlvu3JZmyUSE3ILQ0
Sy3ftANfLh00FGGZ2Z+w3hIE+3Qx5F0EoziHidX8jaMWXPfhkxhoYgNLpMhdnabc
M/DjKNJKisiLq58vefhhKpsvjb83CK0gHJX/Qk9liSSRVdAFEczUrlFmJuHWFsAp
4Oda3xRmMPeBBbJNHwUzcmhMAuyboYNHDKqAy7aDy+s5aJXVHvd6VynWLO7d8PRj
0STTCpgRlfcoLjx0w1BB8RsywsO53Q0k7k4VZCVg1Njv84vjUVulEBuYZU1lVA9X
61bGuQV1OG7/pgURUHkMmP1PWr7MSvX0a8xPQpurAZUfPqHWQrogMGGf5KS0kVuf
rcnz0IL5CSZt+HALDOe0uKU5HTxm0AYgZQ9LG5WUoObQS2rig6B1B12/8t7kvxpg
mD9XfH1/oq1k86QUPhsDx0zlTpWFPVokxmtWDagasZB6XqpO4sAA8q691IpecCxw
3dhtqu2tPJIgxWAODOUT/2HHGpOVC1OZ475uJvKUplrNAb71ibpT9jKM/uDqHtVb
TcY2NEXObQZ0mKbDCPYX2pAKE8dpLpNhqZJB2SzzvdD9vPF3AGWcfWrjfbDlCa3l
vAKps8w3GGJJKe5/ZMOLThFtzUdjSU44zEm1f5C7YCJaB+xUPiIZynmsK76pAa09
nADhYA0JeyT3WTHC9cEpDCVeulXheIKUueEBYj8vNgEEwELgH6sWCwpnzQux0r6o
YUvwMO1s+ciXYHnzZ0S6O9OHvREY9oMdTT8IEBHcsou3xpaDs0AKA/X6OPMhOS5O
+llihzoQEUt/R719tTLtpj9wVtxoaOo/bmG02EXpCG/CvCikdkI6GkUo/ZgmZM1E
wZRiUS5Re+yvWxdq+Y+z+16yj9CyGpVmjp3ZuJRS3ftuCoJBTvQDpF5qFlpMYia7
pnqmiGygpaf8Lc4ycNvwmECYDHLfWtB/arMARwW28bSJeNEpyLPxemx2iIkhWjxA
rTKNoPegTQFnwdi/6b46LUQ0MO2C1TYk4i5SLysHRc56cawRY1ydRhVInEKm/E3J
unp4Y5SyKTg/4jSqePb4u3o+Y/2HKuuqOwL53L3rNALCNGq3ZPoOSWv9osIInwnh
KuJj3Xg9HmnTmqpUZSZLjs+7gMEl3XZ+Hp6uSQ3qsD5uAfiVolHEgNpOYnnlU09t
ykOX0WTgbBrf5fC7h3+DA9sHeORHUP2Hcum0WRsCwE63hDtW8C4G/xNkFTFyl3QD
q66qsMsFcvkWkuw9foHAYDErHuxbWX/Zg7ffVReYqPNl3eITltDolSQShc55nTPV
HKKKVvolyNr1umsFSvZgLhd2y+u6u/Ahxj6bavLL36/kWINj1x3ZJ1QJGHO7bcvs
nFqeyVLosaQ8FdXU53bJ18XExzbVGOpYFpkGvpUg7KGTrRX5JDrsy8qikH9M2nP0
S4TtsLKy0PcxE9bqRGWvCSa6s1FR6SGINDjBiAbz8oR/8ELnGUbx0wx7RzP+Xqve
cFYUWJIQQBkE8bC35ziv3YP5gvO0uEFxAJhdpMqzW5iS1Wnl1O6zhmmAN3uu2C+D
GlpJTHzVoxm0WAnNq0XsuqHD8vqviPekuk4i6P75jTke9I3yaawFeuHuDKFXMEi0
P4/7iRWwH22Lb/gobyANnzANDCocesAdf71zuei4tXqfm0me0KLv0OEGDMKS9Uwc
1C4CYzmw/BKiM4mkoX1vXYrCXZbhetuhwebIO84Dc5r7HIumvtqr8TpO3XlTuJ5K
7KzD7v4A/LQ/naaczEfJN7olfDCcwEM4U94csE8Ry1A3kJV6voyN3T+cyF7KTK1L
mB8tqXNQdEKbOtqlwFBvJY+1Q/v4PJVzTWZvQXWoQbQ19tMwoJhfZl3UL2kEt0uN
wE/0hF/fSWPdLzm4A/+4QrH7/UFcew6M3AEI5yUBeuiW3SewjJdfxHFUrkRqF1l+
atzRpC0ZdS2RU3EUn4JvVQLDCe/QvoRSB1lRu9Yu5tbZV3EW47KmTjloTMmg5zq8
qYE4ctaIqHOybK5Way03HMHjMWkCSRCyw2PmhCqe4gjr/seHl3/Q08Li0tHPUzH3
OjwNIZ6gEZKpITWBCCpBmrLvbf0xq+Y3MAi7pimO9WgTHNEvPmrnOUgtaam6gAsJ
5Hx3fGMje83ccRmDiaPjiujAiKV9uxA87M+Ecfda8lTyK9YeQeSEfjk6AvUhU9IF
S74qGBsbCiUwKnEOKcpinCuaoeeWxtzbPeIDFouUgTxg8yHPrZbVTMJ89mdWt29P
UCtJWbV1yn7f9pl2EQqVsGLgpEagBOvNgKe8KvvF6vrO6Ker68bGgMh2u+Qw76Ja
w2uM1w9wjgez1atJVnsgXHd8+ehuDOdyiuyTaub4WIjJ4/V8r/5iL25PDsfz1u/5
nvuAPeGsakjo/6d6G2a3UYCY4HBshheuU23PPvCYFj7BtWHWc4B9cgD+wOXQV9OY
Ep8tBIXxhg3fEKDAwOH9NEauQ1p0okcuu7sg1HyE42y3L1LxAYG4hycbp6NcLJDw
1CwI8sLoTyvFS5uUPxVpfcKZNiF8kWAJQBPQAUeGDyqAI+Un16S+Nrfe3Gc4ndfu
jjnuXL9Ekck97ZocEYbk79o4JhKLpgyNwgadgLlpCrtLxLJ1QSVD43uv4fIH4VVk
J6eGYd8C18zTKIbC/nkZY2YxQ/MpSwas0jAMajehQ7WeOQFrmtzqHlXQxx1Yg9AN
Cdz37uf/PgUwgi6C6Y8CZnnRjsoWP8qwbs6Z5zFmCb2VOsPyPSuxjfzRcG6lt4BJ
AItmcp972qsijOU0IrWMmqcD5aMryo0nTfiENrUeg53CP81Sfq7WjQGzRiadftlS
UsYm41m2Oyv1vupGi3o7xvoJ5Lm5MJhZg5sDdgvuwe3rOT7i8gK++0AAAdJD4apS
r0WW5CchyS6m+O5x/Kgyxj1zC447CvTkd/TqFZ+uwRrtODFLVB3ioOYaBWU1f2FV
z7bx1eOwJCWHNE5OjRlkzhNKahpMp72aOmJ3IKJmMt7EkFAcV23jhqU1WjLgPBdd
TnG1F6LWa5UMAUKz8L4yqwyfHT7NwwVKC1XfQsBEtUBOA+0Vv/ELuqYOdNMksiX+
cDyZws4B2mldRDtO+p88wYkdTzF5ZXOjiifmma8TqudIwnU0sMahHBDd6CZKAVZk
nflVz015y89NakYGbBesRqRhOhTAKnWDcrCXfY3gvOZ1jQSC8cNuEaLVkfYKelPd
BSKKZdyprI5UoLEMa8Prk8Q4MuR/2LDafI3cojnjbvfuPaeXD64XUQVhPr4w1mP2
m/l332NPQk7Dk2lEZEwmnx58aY8kZqpbGjAd0AzL54FKq+c9nbqneHb1lVV42ZgT
0+GlHg/gTs8X/1hHXw4xJr+D09oIQL1HvmtUXqSJF4xK558omA7lfPDk57R73H7g
/3zNC7KCRvBWKxDL1hc6bfHm3CNbqZRRwqBnKVFdQO8GTx91lanHoDg+42/EGRJR
F2u1QEdu/jFoOc6aAjGVq7NMIwKqSgujACTuIVHhgANwutDaCO7vcbbbIkch9PEk
S4C9W2Gg3WvOEsJnMm2BrGfD4Gbf2owqwEz9j6U7H9AtNYnTmTyijEHlN9eDg45p
EQX8VSmxTNzxpjnsOwQkaevHXCdD+2FlyZl0vorJumtmJdI9YRfcCCsTvoPFB4sj
KVoi6vcTf4K6A4wNKsZns5FME5YTQL5iKCWbN49QAZVCFol6QwNgp6rHQU93z8bX
kDNADFpKTq/7BDboqoqjTjn/oVd3zxAcEUbmzHBVeg8lQeHjNxSI/fvg3kVidj9x
V3iIPoJaMEWeNoUWWKwX7Go4zJ55h2KOnM8EBmqTac3yvpVmZRqhyJBsjV7bjwuM
H8+Lz9ZbaH5R5X+WRx+2ufi8CSKIx/9RHqtZJu+RVdATbP3NlVBVnRBeX5mm0d2x
rENwGF+VRG+V35mRrqiqd3FD7mPLZTBSmKqWcaMBV94XvZGFaDGw1AcHn7urHPIa
KGXHmkuHCu/5rWlcCfuvT4JRY2b+jBpBve4D7YX/lqIhDAiIJqdvqFt6HK1fcpdU
/w71TB/ndPIft59BfJ5OzWQAKypl7503xJN4fFCjXjWjHkUGNwmMpchtGU0l64Y4
VEbExVisrlaJWb5iRx1PzNDwR6fJnAKiudhiea6b7IBHkevXKtkaG7+9BRHtjaf2
Ke+DoarL/6HQR35YnNEctFvD5f7y1h6ZOtOsKaECl6SgRjT/C/+sWR189dXxBTea
TuZ0uC8RfMzm0KWbuXDjvfkU/Ptok3Fw+U+AGPldczS1pm5zRH+yReCkJT2notcF
4r4+ssyLBXJqbU+c+TIDzmnzu59ijtPNfeFnSXASPw/pv0ZnSYeBYJGiwIFY1yus
dsAPEa1R8fqCR7ibd5DkqHhYTjsBHprKIMnnqErGnfUEi2D3oTcBo2jGfvPe+xjT
c1CXTHCkTxSB3PoF+iANhm7oWD3zLf8TyxkVx5Gpd3lMdt1d1q6ppXnPS7VVjYDW
c/C78u3wFZCXr2wnV0qJK9Cn7a3/3EgXpuVE6Pi+twS+fGEG6eLw3Ea4eAKXREBz
8qVsvFrwb8kEkMpCS8TsvS6FTUtuM2/84zK/ki7qcS/k7W+o3YoJCAyOuzOWc5ct
TkCCOqzn4pqFR75wnI/THRuHlkOQ3HJbwWukELy61jx63J42lqV98GPKJAk6bzHP
zimS3DfatKob0pEhfOcjPISOWMJVMsyUjqvRbDWo1FCvLK52eMuzcir9gfpTbsjH
CbRLlovKTY2mU2cBC+DS83/1P2NDqsQyv3Oit+pKnheUgLs/8iGR3QhRg9aVcmux
J0RJdvpyI8NInVxgjBBxowzul9100kEPqIrVYDQ0NLYMV5gvkfKoIrSSlBbGy1gd
4dON65LYAEJ4syU/KVkR1cVXwBkzPXcCOf9SWRDLeqRmvxD7YXWJUAiV2LLKt1A7
K+Vg7j/OjDi3NYo0TFW7pCfBZNq9DnXYhVrvuOScwmxUqPrT9UCaRkXAnSQNd2L4
mISUmB4zYtCHwrE5FpJlaxgJLfP1B65baO7hKhoEMfSCHb2gk9UPI0YOzhiePGxy
nUlb5UOCOV+ortTI65FNv8hpDiVHG3rxdmP6SsPTN2YDuaRp2GLIlvSMOi/Dy1gm
GS1IR+yKNuKhENQezuJZB7ktnfTM1OV4Y0P+7NfEKfUEDZgSdXv+c1wJDfHQU+/p
HbekdjwhuOMtOTSQ02hluf/iKB5TxWQ1KeD9Q/t6uIPN+wuu6DfL90j11YYQrQYr
+WXlxogKfgUWdSAzuXV6o+G19NzVsNfkBLZu/pUkP8SbK7iCWcbdtZaDJzx6auR5
Ail7VmDPjaG/8TAC6EPQ/cq5KNAgUEJbwfiGvyVXO5th2+EVkSGTuqPg+MStMTak
P4a+QLMbybW6q6IzPCRtYFdC4Dtbku/MRNVuoWROCXmu01xNj6ZkvGhcFZc01EMw
hIih6oSt3ceOuye47RV4vaAS2aATNwTvAECC+11WWDUA21jWNQILw2taB3q0Jic2
fXX+JYf2SDfz/NA0zvAU7X7VygXHMSOGcRXC0SPyI2GEx8/ZsFEGnMLbAqDVUw/l
JbrgFmfDZjKxCnq7IciIystjzPx+sI5JpZ4LkaFzgWsLgIvrxajnOPpWgvUOxiXH
z9zBuk2LHp/+kgPU1ts9r+ykE5hFagbUZkxcCHvJXZLwMiiqNbymAACTmmrbeLNq
UQX86tSPnsKWs/2wRYjvtNI29MvOGubMMM7fnVoXfKp2DmTRZBs7Wg5J5cLGUlS8
X9zNOH/NB2Yg7IybyzD21F34ZbM8WqmsJjxFSiEmNSU/SNd3LGzVUQJsqpslPler
CkmfEPULnwdQF9mehmQDG8MGmru6x/uxnBDlGy8x1Mm9Q6pFM05ZG/TOXo1naZ2X
kFQZ2RienNWJ+BLQwyX2TyrndvogorSM39NCiEwZpYEeKht8NlDUvc378pjzuy+w
HV9sbXWnL1OtX7QgP17zsZq8Se66DsG1byk+ms2jOYswHJD493UwsUYXuewZuP7Q
BrLQdoBRyYplJhpxEhVCWjAP0lvTl0cUR0xjSSbq7AZLFE4kBPrCreypePCVN/zw
j1BAZb9KrrouayM4e27m77BeNcW53XkfGmZTNF4W73NQ/Jf2LAaQlXP5FhYnsLjg
Hcr1sO1yZ4iKAliDE6bhGvVoLbklnH2BLYY5ddCTWUL75A528TdXNA1uF1lZX2nY
ZAgRag//aGB5HBxh22sL41P7aeZUgGKfbIKzOXu3qIjmBR9KmkPXTSI2q0DmCxpf
dL3RQ+VosC2n1/ZKRvEDkd44dkMdt0TtMJjNhkcPE9t3MF2iDshr9g3x6fhfktni
81PhQce5PQYu3TleQTuEdwooyvR2hXFieNdr1yivvXDRvSwFXsFyTF6T207WR45p
QfgfY0AsBJab9BpZ6e0Op8PEuWX3O2s8IeqHzTx/mbnZAL586E/20pWgqeRWGUAW
7RRUbm/1Tpa5LRROBuLdR3j85+mpisPvURwJXr5PmUY32lqnTQQ7U12JgqUI91lL
uq8VIh9BRehhFldaNHEuVdKU30qngFee1GGk3IR0jShUwNfID5ET5JrKajBxn7cs
XCXqogCwHQOsyMDcBowy4fzH55qJ7EckaLKyvL5aTAy0ZiyLX6rB5KP6S201z/pw
6xzlkwQ8d8rxIz1NaM0UTk4Y0kfRiC615k5iDqGGs50hicOXBwKaZxs3LhcmuzgU
s7IdanN2zjO3V9/ti+hRDy2Y71I/gNysWQPG1acN3GExf15NatkpfFa9NZYYxCiy
T/zub3/LBV+5+xw+7CEsfuIrAYFRyMKrDX+lXtIyjV2NWSIHvtzUl+Kv0/1oL+Qe
R71J59xE+gOTzB8aCVZZghMx8b2tzNvtH4pXpVo3rREcirNjD56Z3eHyiowOkaDQ
8JQk7Gqkf4bCjmhVhE1ND7BUrYSUQ36pwTJrNdMMudrph7N9npvLpG+gY96h7O2o
qW+pIT9RdlvQvZqp8qlPmzs9EPw5YjQD4v8PgX1iqAKiaVPnOl/qqF1GmnAWxFmm
a9mTFCJzYUUrTsbfpktUsxf6nnUhdFjtBLElgTCATGtSZ5DOEzxftBu83gyYXbGo
XQjRflbxA2CMk0tuvvfjkuQ6enqW2QO9xq2mRs0E/NZV7TSl4aGl7lDF8KOWd2cD
MWvqDd29xnPqFvLKDpZetNjdYGPlzfzTQwGwkFP0ZdPsuA33c+kI3NzAwhA3UXkG
Z5NsGltUQ3k+WzHLt4nkiVLZ1Sd1jHC1Qpnfp+tAleyRQ4FINmcf/enUrOGYilrS
ziyXMu6pj9L3Y0XbDoPDHEe0syC2V5oPUow6eMnyg6naBkyFKw7NDcEl5UXgjx5V
oy/Yl0nANjNQdtBacJO+x/vQvxSA0SCBQEzy4Jv43tykJmn9vi7zk8/GTueu5hTv
mQFNIrKlXj4ylePTW8CYmSUFSgqNDmjrAKCNxeSxLJ/NbZvvMpcbL1nsu5byE0bh
jNEUeHFvJvIGvS6M22QNlG/eB/PdW/v+iju8YGPV5GZXWIh1EQ41+mtOBFUZjxqH
5YyJ6eeGDtA8yTeFtqdIHorBuzdzloH14xY0v3zfgnPUBctj0UmCO1josodxn1sB
P8bV11LrucILw8AAkFt8wQoeoc9TFfDcPtYvM20Hi8PGWGykhDEHu9KKHlOg4wHM
+EGc2f70vB6OZn6B6V8cqGa8ZC1o7pL+ZPHYrxbMH15mZ1UTP7+lNwC/nyluWEaH
tJxHzQbeJ6jf2EW6d1XWFENFbs1IIcRQdDHvsiU+8zqhY2H/NhcqQRAyawAjujea
80t1CTd3MwXCmOs9kF5ndtZiJsYUj3q5l4TApy3k/yi1sep54UKiKVE31r+nkmhc
p6t/EMtIsNU8hLmVE7yDmZu6kcSRUEfGMKr2gBxK7rdYv2ZbO9xnePc6WPU98YXs
JYwK1pOOSXFcugnAWJSmymvzQqC1ksVM3zF/ZIDZL5QcEPcyyy5bnl+WwzK4xZJ+
lCW1eVgRJkamKyVMFX/535rQQghu6O99eJlr4nBz3aULfdBz7vQUySEzYXJuKMYv
TquF4wLE6boRFmhJ7QZuFbxbLQj5iUrVTwFkD5ouNOajBJGPyu8QZaVYTZZqEEli
DnUOL7jNkzSW3pw6fszrYxSjIbGbXfa8gZHOlXydcaRa1wSDb1VNYx4o3rNx3QX6
YmZe/faHsaSM/ptihrNf/cVuoBcLbtcrAKwYoAjyIeZO9ZmYs9VDiWr1zDVrNmSR
FqHaxqE9V/gS0Z2rsQ6wM1P7LsXvOFm1MSXtICYnRBvRpwUGSMHbu4pxMjXNkSsv
Wp08ZjO/pJRRCWeC4neYRPXO6gPMEHMaJ7Y54lKnhhPfkWzP0jLduD8sKhAgJ/oq
uTCJ4m4sK5HBCwXa5UvJH0rhDuE90WMsAnDm8PLyp3I2I/aoySIVuxc6Hzni6n9O
4umhqgOGOgzyb8GZ/1Xz4PkOwDL3FvekSS4LaU85/D4uUqEVv6Jqz5JV8tt+PLUX
i9dRx2ISUVanHqNLFp550ELiMf/STGExsqJuOtsUCcUnqI7zYBHHwODY2DVq0wcT
fSaDalsXv2UnMOJOT/dYzkkQSaNS2KoHT5JKYtXPJ7vI3K7/q2D7H0TqvZumI7J6
7v3Wy7VVRm6YdlSRZc3s+GUrzxvVkRMyZ1XZanrb8majdQ11kK5bLoUKgXJKhPrL
8pzV/Cvba5q2iV4DzIemm0cPNb9E1r3xLBYrm7lF3co7mQjEeTbgo94BiBwXSsyf
18KnmBMEogwnFe/1XjWC55JKL85gbFypI/TAgHW3DbSOCeLY+VQz+9iTOtrYCCo0
wdFFShS9m+zFrQnAqW0U9Jf/FY+5zsJz5PEFefi7U62dupfayhiLSUAkGaabYrbI
iA+gC2Hp3nqeGKCXM0wuX5ggX8GaaGcKHjfiL4IQqpjHHXSf+CrnWzJuOMxD5mEO
2RbMqN1FmZ8F5VqtptELqFmcYilU1gLr26pZbi4Ps7a8lEq2yxdVL1e85g4w7Etq
uryThZMmNzDyDYXXOXykEZST9LYqp3AHFUiThBW0V8d0Au3fMbhdMAv7WfIhU/t9
Sr3N9x7loM/e67rfDx4utnU+d0x9VnjUUxcq61pVJPji6S/uC9wKs14w+Zfr31pW
jfvmecuEuRxD23bW8fvfiFH5ggoiGy9BCi+JLGAGnn+BkqE3vV0Pl6ABr44KxTqy
b44OtpLXx+Ou0tLjO1Kyfbj3tkaNsaM+5zjBcGyZtrkRDNM7UGRDHzM6tl5fJ2n3
TgbX6YXOwuJO749/u1caS3pUTyXjh/XY+dLnCzWa4lfAp/IB/ocGCB8XgbP+Cwzv
fuLA8q57SWl8Xd45zNAtGRrlrUh4mvYXXHeWI1hPD0/kS+g1asEvex27dUY9j/8O
BW3FOvjBggaffN9K9/Xgi+0XAoc6JVYBw/OOouPIlTSMrANMte0xfjO1/TKhLaxw
LzTH74/FZSzKPAxQjZsuOYhCQtu0HO+zvXvZ6nPaz+/tyMwBMqySNiI8dQbWWQ5R
SxBH/l6OVMa/IWz5W5y/2r15/yFUJdkedZAkp47S5jS29tTkgAt4nWGuQWJsP2uQ
JYmzZ6zjYuGLdafwtZ6okdNMQZm1/blG/LOp87KDtj9TcGNLczeDrSHruwRcDh6q
kZZvqBzBgY9iDmYvUto9YMlgrv+14vcEbAvOpEz0LLRUxWdeIeceYlnwOGWXcJLJ
NVGDKZWW2OcMJp3UVTio+9TugT7szpqu2o20f8UrdWOyFfg8+4yYjISBv+lTklM9
Hap+tvqcmZaKKsCoogX+FbJP2gUjgkqoNqLI03ycLuv6gATN0QTtKaLrKGQRV+8Y
0WZNnT9Swg8hk5g3z6O/CcMWsnPMttj1oIfUvlyM+GUp6qY6xq7jHbVtnR0WB6sT
CotJCPZlWGUIFOIujJdApuqlyvE6cvY0n0SoypiRGjJeOsSSqFv4uzWcKquYQ0yT
cVI+NGZfUCqmPrd4afpMsnwH2zYk3ae9yfAcfcW8dNkLhc6JA1SOYc6RbNicx/yi
UGjiH+a3WjyvHaWDrm929SRdYBd/OmmP2aIrBGO8uMt5sP2Cm+xv03JaVGFiJ7tZ
YBggZPe9NDy+qk+ODLmrLYNpESUWckLHAF9Td4yRAuhJbajG+pyadt2oiOmJIoqS
V9WMFWN5fOAtcI5TfiBxSotuTGRsPDDC7V9KgIHfkyp0zl6d4cfD1Vryi7ZrCh8M
t1K2YdPGVCvcbXLrmHypSvdtYRucLnFyFN2jFcQaO5Ll9jvGTiuu/dnL9TL7FNv5
8Ue9J2LOI6wQkzYc7ia0xt/Bx3UbEGMA89qmNePzF2w6JwXQpIqwXuvYSVr/L+Iy
S65qjrA8lFGs01bYZNDIY+bpcm5Qx03WvnaEigrv5pHgVPKkNmhYw+H4eQPe8oJZ
GM5o5GfOOplMNl2qO6uAcGY5GLyobTFrdF0ZfvWNr0bNFysE5YOU7iiJ6QUYtmp3
gWS2QhjLXWEVBPgaxTZPQT6cgVtso5nv7pQqlQ8KV5lY7yaL0uloxEEnh28EHqyU
4CA+PnfpzauKMFUctg9j+Xj9JVUtVhSW3lowZezE8MfLoZheC5EzEOqX5D21bqJX
ZbYcy3vtHiOXsHSTM0iw4yrXm/wQkxtNJRBLJP75NAlWKQbq24x/zSjliDvmBuz+
5huApEDk0MxpmuKEPQEY5K/F6jKwlQ7FDBtlLkIuYLJ4shRqTSlI1Xpf/oL+m1aj
ovLKO3MeHjlnnj6HLYVwOPmLld22MdED1h7e1Zu5/tjX+qRlDfZI1Kk7Zd0wwgKt
ntpoJAUrBXMGTNRtnwTwhm8HZy4qd/IlmAA/GTbQj6PiDnjfyCy/lfeHfntaIDoc
ee4qTII2/d+3x/GGlz53651IQrpBwMRrETVSZwZQz0E8LFkE9HqpSPHNRQ/TBK41
6uBZzGhFOFw8cENIG+7hWGEAz7JecFewECAl+nI8hThpvflJXnP56Unba6/wSMmT
2jLvkvJ4/I7SGUBPrRDUWpU2Fe3eKmBGYN98LJWCvkrvzLLtmiys1CSBbTL0kHFH
0QdRZBKO+aqgI4dCHdkSSRnwNXcU0tJ4EUuXuNKseG9GjwMAk3FeXrdZnDO2WDwM
pNLoK8MkOL8Bxn7QyQ9UrTD3TyARxmG2qs+wURSYD93Fiid1jh2gAi5QKp4k5xvG
42ftaeHQ/2ypRxK/fasoEk4uKTNfJMmCfE+elLIHivhM1tIc52fpIrOR0hYlCar4
SAWMAVy9e/m2n2PolqoP5Exe5k3QUAjh/xyN+6sSF2q6OhjTmTa3pyV5HncoSvFw
BnUV708wFjp4q6EJIPgf5pi03fo9HI3mZY57104x1imMYqjRoT6pnZDOB861kKWH
n/d1YyPp2WZVu50WxukDfd7awKxe0FWz2izOvSjjCl8qO8ZcrwDBQ97OAD9ONIdd
cFmlpacQhfcjAbhPl/pl3b48t+nEexYaAIfUWax2AyFuh2n/dc19+6XMr6hxaMKL
3rWHfnVRLgb3cJXA3ZMB0xMEUAOt8cRpBt8Fhl1RulSkMwhbL03Lg6rCKwl2hAUK
U+CSuys4ImTIvSDpIU8YO1N9TZ5IXw3fxsUMDLIWAgKjHXMAo+ogyQU6LdDzTiRf
AVsxqy2/W8pB94Z6YpW2lKt0OOjVucR5ZnlDp1TYQTdh3mBZ60+DDl7/X+2t2KND
LM2P4a85FgfFx8YcczHwXY+4bceXUhJbaT/KATDuvmmW0CSU94vuiPvOa3+vzpi/
HObDxYMR+AttolYw37QA0y63w3GGHpIcUCwxivd34eE5bdU6m+KdzgYKPx3pu5kr
ns/r13IFh8/0InuSLPM+UP19s0l1/xNN9C4aZxd5orMIr+RHUmlCDRnGDDwCQPbg
BkVLdWvMf/GbM5PTeA+ru4ka8Cj68ytk5afKHF0MWPQWyYijAS1YX/TYMk1x3NKJ
fLKj4KOfxdocw35zjgTdBVjndd6vfgyF2KzgFIkq0UQ5Nuzuz7iiD6gZCsd75d8N
r1rztr6NvtS4aKPkQXfAm4P0P3ekq/fggwBYyWYhHjjFUn8y9eihJlDqrsM4+H8F
Q17Io8dqcV+0ZOPREgcGfdPg8x+jjoVoMYb0ux3p3bBXkHPfwfvThAr1daKGoGnv
Hycywb8aWwhWSNiJpHduB1NPEk3bMs3kD8+rWn1P/Vq/L7xCNDAHL6ldQhQWwBo/
wHWaywas/Za1vI4IqnDrf4MTZEJPIkk+qgvj6Wdziy4tRx0k7j7Iwsl6QQ7X4aBH
AxuhA7PFTLenZjYYqDm1Q+tJGEQeCN4e9n6+wMfhKVsGijXVXrosNLfQm8mSbsvF
OYIW79LLz9T9MH3jFTVrUSFs2XIs5ZIfUThVxTNzo1xHjxPXa7yBdUvJ0kkbsLS4
1LLzvxe0/DRFzUMZ9lmc34c+V6KOieMYWezJvxi/IYrj14g4jordrMIZNSPJeod5
5gSFf+qFFrjHXRkYbZdwLEdD4ZfYhlc7axhZsJxWCuQ6QLctjnwIupummnphsAf1
1j6gOaa4lSCVFtDiXBa4nKgN4fqTybfyFi6kE4kvLRgylikCygppXeVjpBIwb4FX
wDOWR5CviKrSrWPShD7HCt329nXcTCsaaWqFj/ELLVaBOpjXNGjr46K3+z+74xeL
oPcbTQv/f7f2HnupIouWYrnZ3bdEAXPXiEIRHtSNdbGURLhy0KIX1GDjIf3WH+yd
CJu0UguRJub22z8jbUm4/E6gHBDiPZuVqqQihImUBswZw4T10IcfapRUNt3f1e9K
fwYy9HWE4PY+CygI1+GMuOG6nL69OieT9ZED+o6TjdiZvhXvonByY5Cx9/5CzxXQ
4/P3SLlmvdqiKojKHBTqXkgXOBs6C6iPkcSKUd3R9piuAWc4C5BhXLstcXSMuD9z
y2VP2fqjgHsgp6Tu4ZENaxExsVGCIhaXEraTjTs+p/I1Xn9km4RTQPY4aatFwzO1
xsH3TNOS8PFZlHL90hxfE9NyOVwep97KyAbUr4BW7eVZ1Ff9yEdFQIobdl50Hty9
fVJi7DXS/aPVGt3Tmqq0Iwib9YeUGbfZfvvULQEVNuDWsN+wWOZP/LiFHFvVvqSi
QF+dPprFBvhjAgcBbHSEmZ1ip/PFAJgIFESrw+EMrBNGBkTRcMW4FZ5+VrZU3ewD
Q6YJ9TlmLWr2MFa6HQ5p0N6GCdTzhPIIpRqdZIePQ7LJ+LmkAtJQO6yKYZbm4Os4
mjZoR62kdlNsheiZ1l3JNejP6an3rXzrTP0enfuBghjwzYdI5y+vfXqGvUW8lJP7
HTz01bvhlGGMxX3ker9cdTGRaHAksvEtG1Yh4Ttb2cZHSFLWcz+hkMVLV99kJlnP
x5KWCFU5RarMZ/o4zM6ks2nAX6hZ3O3WPkvR1dNZT6Jfw/8RwsxZRRJ8EoDt920w
ZduUGYOPKjCwX1PDnhDXljImQM/6uDRd/VLwP7zDPXzeLHD2RB1b3hGiX5lX3tYW
nBAeg3RmVboBl+fLujnr3kzichxa3k4/rS26iT9lAsJEc2Jsh5OWn+ohiiHllDJP
KnC9boQ6UOxL9YdvRSDTW5YAJp1S+FOmHc4Kb0kjSdR/FgENNtsJHP6Ti0aKCwlz
Qx+HpGdDhwMHLpwLTNPr8XOqUGneXZv/w9+lVYdqY06QcS02fpKctU7AOMFSPes0
+QMUCWzNZtrC3WylHuUZUuQSdB+P79ysUlJBA52B3gKPqQKEzMvJR4pZP/YZQtDq
9S9BZq5GJzjjN4S1egwApSRqh4RralJ/Fdd98kiQDF609js+a4dxeY2nUt5t6Vbt
wEXxMloOlTMOxKzXGa8G6gFGCxQfGS/6q6Lr39Hm8vH0nYwoTWofoDHtSsL334V5
NiOsB1qolS2EjsNeXADhQGhMchUEqCA8KooX2A0T0hTXz9IVJ4cbg0efN6wu4Xcz
E9zbVV3iV52Nv+phHOIXa/snY5WoSAsDcrQEmWZfzxohmMRWuzyJ8H8qJDfkSwH/
ZM6hdbg7UOM6369HG9zLbYbp24RGRYvV5LAOOXLuEMezhPm3vi9TVCrlL08VH3dk
2u7+rDbrEtOLraBiJngOdkpNBHp/B5jvpNR69t6WG2EeqsLuRK6M+5zDqVuGk8pZ
VG/PhnnB0bnTeqi+jqjm0zjRhAYjmbMpl/rzDE4q3qcbWCLoWtoWouuiwrRrr0sL
W3N9IE1g3CBh2Yor+6NzaMDIe0H5pI/NozShNGVyV4PUJpZ809hOoyD3szph/pID
WTa4OjRSpFTbabpgiGG/EFjoRlR6Z/UGboKmwWmUJ6sBW2r94SoTjHCrNE7QVZVr
dspnXkBCk3a2bRkWYLlDV1nCQiMOMCa5aXHntB49X5hl/waN83wa1stY5wrf+x/5
WsF2r6Xs9Ht7j7HfvsWDoQkkBR9qX6m6BJi/QyoOBtmq0EzayzMGhQ7nWbzy4r9e
UCqe7pBab3HeQOs6q+k83Hm+B5JcTpskyW14FfzyOxryOUtC8IwH8T/TAKKgcrVo
0rRaGGQ7tzGVXebilzo8QZqym0jrnxWFohMPLXmkeQIQOgG3ADvSAD8DhUPHnsbj
hIfA2hPqVvgqwXWvA+s8CtUGDyGPATGyYwklT70qnyAxGoHjwu743ujgmBSX0XL3
7qQFnlZ2AkDcqu7c5D5M6SZmuClhbO5BAreZ33tG+bV9f9VYTXEvyiQicn62KOTd
aZFOtBxzmWAgYhgyyp4A88HHXkDWHTDOH6aewyQfyUM8IFC2esoQV7qtgDkZCfYn
MXgFHxQPmKKm5IFhHvzFxY/TxKMRkzsSSKvuMSyDcE6Cvp6fNtumJjJKrqOHHhCR
zq6uOQet32OPQ7zq2LbUXm6Td6aWqPIquLPVJdHcDhDgGUiwsvJLbPod96+5eDPb
GGiVXGk61/TlQrt2j6GofK0ISG8H4vcbIRgBUag20I1Z4JNhw2eOUISDuBRcYAxc
0Zr50BMRSqXjhSSg7qjzzf7+Pdoqi0GHz5Yq0wuZQDz7cFBq37ZZkl6gPgqb4z3L
7oNZaRqf71SHr3933DbVwbwFEkcklpcCLlpHnWLGgFfq2CIfwqusbO0oUM8GonA+
z+EOV3ywMywxWbmoLuBN3Oa2LgPmjdmz2ZaEf11zsRL1JAFeccl1wnOL9g9As01I
LkkCVpzONo5KyAbFPkVXPL+6KeDjOKs9Hlra7RPrxPncrwWmk/T1rMCnNH1ba6nY
mdSb/O1/7op6kqWYPJgY80ZpP6TBxdy5eMSxb2cJ0H4wJLDml3Ym7yCHwGsJecQd
MgD504pE2J3Pb9hJeoHW3pYrl8qVCdw3twY0YTJ3sQixq4hM3Y9TiJt938HueD9u
dEmer3H/an0TiWVff4UPmcYZs1VlGHtHoHFUGqfGtQsIT9FY7RNfsxxtRsBw1IHi
dz8JR4xwBszK+IBorgTFWPZJ6KdeORRLE14tBRAYSJpMBUU0vuHlsjrDdheYRlXM
zFRfLpaih+v7jNgzWCXOWTbzqInhHhuwBMXdhRtcTpORQt8aOzkaNqnAMQd7H9Rc
kx7fuMPOPbHMicUSvhwLjNRfoposUA5tnD/XztPHMBWgQGdNM1lllwdjn2Ry2Us+
tCKqNTVIoy7BoEt5aeduqctFkxNFnuFrOYQsu2u2bdGe5xKlUQGOqGYhrmQrhboO
15B5+fj5YvEv+PRY7ND8zBh2HH4UN/tZzu6g1xNBtzt6qYq9zKR0jaqvV7ZiQprG
LlqadfAdoshea8p6fya7hgM35DvNRGkGVJF6QHQkSdbBZWF2Fx5xr08SfhCLKgH2
NJ0ACsUFSoDDcRy0iOySsPS5MwYIjye3CTB0R8F+SW6IbmBZqyZKMODHGxMojHE5
+34/U3WjFE15zZ2QH5NpLSLlzU3P8m/faYEUu+AlqbfqdapDzKW6T950xB40sVW4
TZwwb3RS7SlLWWiy6qcdgR4WnmKMm7URkgPKKRhKzLLcnVOczfli/ATQahIl0lNw
oWNy+nWLeeTWdXVl8GlhytFfD8cBulrh2hoJ7J/A/Oq4xSXQLF2zdWj+l/4qYedC
yuq4ovJiMHSoC86aa1c2zcId6N/USPUpdggTl8k1F1IyeHPHkP9z/TrY9Nw1HQuu
O6d8vlhen1v/DeimoDU9XI6tX8lTRW9Gfy9OAn/t+6OvTaO0Hlkj0QPzVVBsrTNx
soSGYGAposONXvQKHmcLTUGkF/Qx/oUHTRA5uf9abb+Q4bIRasgfTNHBCum3wtDU
1k+unplk2R1NoxzxConXZmps8XnQrDgMSU4EpTccFo8VTwtxtA9AThIrowW9SaNs
9R9F78REgcgxTmjO7/dHuq3kGi9kUFcxTeIRBOQzig0EGUNvEyiCH94ZHZlJrvnC
8InChaWWcTkJvosBKgRlgeuBakJ+uFno+3qPM8IdsfQT6ctGz9QMzuMmSg7WyYwL
MRLu3eBiObQreCsEnGAD2FmTTZAzyRMrkqN6Hzbwo0us1iPsOhdcNpCkGR5V0OwL
glq4QONyXZNQu5+gtX58tVzEXErUlLYgMkycRkPTc7vfWx3AQ99tadOae2Q373cV
ZmblVjvTYnBP3lw7OJywPZt7R4yTPERUoMvYCuN8UucStU8CzkOoLVyrcvDuJgqs
IztZIOhKPlen27D1hjR77+rbfQrYh9hMeajJxb2DVvebyyFY0lkalXWPYA9YuMjl
WogsesTvYMVvHlG3tJ9OG0kXj4h4xwHt9teYvF7dBhG9ldvbSP9Aih4fFKhooPwV
r6mWvRenP2KipH2yhKp1H/zlSoZxV3p6LRkebk5Z7SF9uvDm0r7TuWZwVDmwY3BU
37Pu7xVqwq4FKhklM2qH8tj0TGy8dX9Fg0PORuoZ8b0c9ivFo8zjKw6IYI7Y7vqO
wfw5jN/V01E35trI25ctVXj5Br85TAWFPuuVIadaOjD3CThBFf8YGWkanmiqk9xu
yntT/qJvJlUxhZjNiVn4Wk8Ubx18UrfWO2nYLRyaYW8v1t4V6cT2BQYeefoiIbk5
nDvjXXdESffmzZrnv/QjtQ7V/B0BvLVT2TXLOqdFesojaNbO5Qs+4Y5iZ3baNOBd
0k6rUTxizwKEgR/GmA3nytMfeUfH8DHrpA+Q/STbg3qc/0ezrpl25nbCCuTBE1OZ
k8ehVoTZsZfGYyjcvTLMTUhnq6rERn4fwAq99JlaqpOMt4t0vILk0PgvV142vgef
G/KaFateOaGn3Em8cHRpVNEuMLhZhruoYVvVK1uL0Ar9KhGxl7c7OjiKbhxGoXGW
YuU++VI+MxfJXpCc+Vl19ARxM1xLo0r4F8kVvKdHfltCdhYaz+oJ13qcysJJSHyz
8u1UtDJg8XpLRBhJ2n2ia0uBLr+AOFwtLKKQmxN80eZyLNeaE5B4YvenITX65YFm
mLgULd36f5tqdYP/gBMJgKm1WncVprErccZh8h5Tc5tiXaGgC1lTwRchuUNGtrj6
YG6PLPX3yc2uJJiMza2r7ILzuQOyu30Aj0SiIohUfBH9f75Lww5TKquh/MPalqgt
QE2v2POZdqtRCxY71dSyk4p7146Ul5zplzPys+SbV9kWx0jr6NN4lEGEdnElwnKx
ZlinVNJEHJSPTP4+vBxFcpBFxXx9sKqedOIROnUF/r8yL3csC8p3T/7+yp3AQnRI
rpSZBukY44lcncG3sAseyQU/XGpO7eVV9LRN6bO94yliaqIR+u34J4cTvdl759qY
wXWsueZtussObbz4sJtaK7v4FrOfaXsIGZVPWe9u0GKqbEvRSXrfU1Ffbt543Zsf
3hiFlbalpjGGPUe5LjIEY4bhCqyucO2EdzcGUkHGNXwW1MYrj0hVu/j47pnC1+pR
XJp/EpnxWKw66SHuIdjou3VivkSBpywC5xgVZ0sKzB29QbAVoVYzPIUcvAiJae2n
vD3DCU69oBKLDFjmyx7lx+E8jPU1LRlTsuG2tixxbf/C3aaXPIZkJE48OSPjzlkI
/7JZIYDzpERFN+mIsWg6O9uzIMhbfNzRkMNj/yGPquyzPmVLiIlMsjc16u3JIAlk
E1NfNnOLxd+3LQ0E0iwsgdKPF51BhzpC/OwbdI5v6B4gJxe95JFfbaas/pDOR8WA
qetvSebfPbQrRj9N6d7oEIuMiOLLnnzZQCu17puSbZkQtzR2y/RjmspoGvn2IzwF
nnibA/0S6ELo/UeZhGYujBADecLKfpJ4TJHUeideqL2/Xfi+iMCbB7RbQKq2vv+s
zNNvu0cIcsjOil4F3bnLKGBu2eMWo/90vs1EtYiKPLt6kluPovxUKBfCy+p37qJf
afQCdMaltNQujjGmQCo6Hb652m4H5vPWdtjTkdHLo6WUPqPOwR+WSwM5f+v+DU/4
FLsiph9b+JKIGT+ZBeCcBcWnTfDBlwmmzy9LTG6zVpvXqwnpxVycvbLKfDJ2F6YK
NEcgU7aLAewfz3oRhoy/J1uzTRDwaQgDKUYJWsQx8T4JYLg3aEDElC0JxxtkzMxo
7ZWjzh9F+d/jSrZg4w4J4AXkXeMT6zuHvWe6+41W6g5YXHrncHCSnRjNh71LiK8Y
KdQ7rg9Avqno9UIKWzq3EECBL+dKhAPw1YoR5Ll4mBBQFibxyvWN322SPwj2vD70
QY3mMV/tOpsM6h8s48Pptio2W5MlalEuqgi9IC9wOeAxJwUuf0azfCAxwtDVs2nz
EodgvSl+twEASqyy+WJtazvpcz9NRfN14ay6EHGxg9Nld127wYSOnprLwMr03cs/
X3BBxp3rwM97CRYsxZe2x7Qn7TOsfCF8cy/xAJnCqGrx92VHNTta42Y1JyQn7rEz
OXU4VXTFS+EqbqcAgBouAxM8lVhEaXPRD1o1Bx+oFF9okkWRrdz9hSeTXd/ln1f/
IpFxEwZotwYNSvKbJrrATfp6q2CcMZLdOoIqJvng1jqLm0Pa6aSWWgurSUmpg5wd
82D87COaQurQLrYYBZ7k1kOtx6nKXtcVjo+lt7Vx1jAJ44TxMaUskBJpwa55zYcf
PM8iWqPD/96Gw/2+3WgpQR/O9eP16ReAYZWYVdOWN2uAb5k6i3hWUltXAjakqEDB
TTlKst119Zouy1gDhFXmdxA3lqfqNrvrk3bISqawPJtp+NyyUiCOZFH0Xon0NmFO
7LoznTYw5BVY7veZyl0vTIj1wwQ0yl5XmKYln2g03djgkUEAh3GQYxRcxuRnmuXa
8g4Z59xEj6MVjltOx4+BjmLRoUQEX+ifX0FLIGibmAEuQ6WvxJ/jnY3WLRCTTny/
9qw2/dwa1kPRLIZGX1+IywSIdNk4maE12BNtU9+sylfBBUTBH/ZeowkyygBOX0eR
ueUvCLz1NxbeE2PC3cXYp+dv79yQydZJBhTH2pIvCJcYiv0GCAouepLenHks5VxS
zoIMxPQ/ARMuq6JyVrh95Xywm8F7T8wp+68rnDv6xalbZ23FnZJgXJDc8tnjGe+Z
rBKJnZD4WPGerJIrEzWFI9xuw72ypXZ9iHTvOluvP9JILT4reQs9S8wWkHfxbkCK
KmWOocn5vAYX1GHSoipPjo9+VXo14nAbq5Eae1wfKkN1bPIH+eY+oUUhn156jtN7
2J1yZMyhHun8O3ysrE/l7LY2hu7tUHcj3WMbqt16OQkHxFYnc+nCRpuSeKCWeRQ5
4apLntrBWTIsrY70/Z5wp0W1WiP5fgt0vJBc4DGVaYGt6xPzaZRPaDTFdFeWYhnd
38mznKLsK+YTVcE8UFg12R+dP8SCbBuiyTgQGcBRQzd84xjk33Kk/67ftbOzl/rW
AXDfh3DxrVC3qQv1eiq+c+KaKx9K7EN2WuCiWLmVtS45sa4VZMcE8qXJ/s3bKErt
yj90YZe3zpIQo39oUvNVjOmgqfNVXA1ddL9WVnpnL4wnCBfYC1M4wf8B7GDlDh3a
qdRFyQ5l1txGUCle+Z1FJgZPOABFTFrOD03lsdnEZYDu2FWLuWR4sOjI4CGrHXt1
IbAfilknATrlryCk20ZRxVSn+KDqcChv8RWy9HlH+g+vfaRzZ+rir+zRuytuOz/+
WsSuYi6rLA2kC9b0SB9mjU9utf2OXToy4lQREky+P1Kys48P4rnrAgpgT0IqhNsy
s6ncJKcssmIExrRlGFxrU+oPZTO0mP8MSr4E9juSs5x6+PTbPMRel+u/0GlJS6uL
UjXoE8D+Wjrror2YWlxjnz2v1e3jlIpEarmvg380z+AZgid65/j2degqs6p86ayj
0bTxuAb2LLs9QSgXfkofCCzd1Ml3WuKMYc4TRlRUA2ebmTkFRdu6sVaGEQ6zNnD2
EtT5luhMAt3FEe+ZmoAvcjlg9531aYYcH8pMV3vQZF6l3uXTpazI0hyZEo1KARZz
vpoHEz2kHpbKy/ug7q0F9joDax3mw265rrxVu7mV527tIkKDFX0Z1KtTHUW90HhY
THy4KIMxPJVUJl1LzKvEucRbmsyW/6geYC3ITEyASQ63X/+Bf9xEk5LKTsZua0i7
WBSa65H1H/g2y5RWQt5pJvXFkyWft5x0gkX4alCfbHWW2/SiE/q4hZ3krap6javf
fj/xcclXnfwGy5hHll4MqX+cxU3i54D3LPIRZh9hVbaxVNQV5clbzF315Ej8qKsF
5LI/D7p/VewEsaHKVQTlD2VhwLEzIB5t1KR/qjxuP9KbY6YYkm6hgOCxkiy6OnXp
EvrItKFZfMG+sP+hwDh4JGCOJP7Ubv+6AIUSQO+hsNlz0GAQAinUsD8Pi5InC421
cCECJ6nI6P6dS9dLU2/zO8l4gmaZzp+5cBJhZG4wkHB9E7Fy064HPJZWv6M/UdcU
Tp/cmvsb/r8aLvkeCamrrCVz5eTaCCYnn3USAUXVkWhspHogcgf3vE/jy24lAzYH
dOvNnGtkLbVoDIw8O9OQ0ffK2fHHi0l/2daKDQ5Zsz/6CfCLBptk2KYpM12zZzw4
fsShr/rJvU5HeX0Ltlnu5NwAepdphCnrIYXzmyGCoq4Hh7q/Xvv8sFrV0MiH0MaP
Nk2m/GvzlP1hFhqRqSvYnQf/zbgaOH0msIUGQtxLtZgXm/rAlX9FdbFmdyRUdf2q
iYe351I/y9DATe48YyRdVDkTbfpmm8MJU6hgSkg8dPe8t7I9ATPOrSXRTAo+sZ4o
zHbd/wGW6IfTZS3ntRX7MoW/1rTlmd9kTEbIg6V9hezZrDBwI8kPRefI1rb57AoH
E3heKEjvFx2g8Eq5QsFiTHC7Tbg2U4Ki0AACemMUNAaROEcm215apx0PK44IrExs
b5GiSvkB0cm4gzuIEKM6qiEhv8gUgaOlo33Ue9ZO2XIyeXp+4ONqDtBy0v3GvJ9O
v0msDMo4PTpcFFtkOUmaOLdB7SYHiuWqtfOfwXgOq+KC3Xx36ddHrGl3AbpNUFz7
JnnMmnNPVWGOaa49Iw5nXXBe3WBn4tN3dHmFnkQXYxn9Bv4lUMeuMyMfmv4OI56F
tuXGIqPrjJqaGNMHhBdswTDDFNTMelUnt2jJeDIGjzZ2TliYmbCE0rfojmYPv8eY
zPN3StL+S67v6TVQfZqtRzrpD3srlRv6Bxkd0cjTv0sYHsGAePHtftMtK0gDaTGF
AJmZXBENy0d9OohQ8jpwd2pgDfnllIAoDP/C1w0uJSIOeNGbwoYrrEXli3Kj5OU4
c7nTbKxt9lbQKKM6706eXE91doFvNbsRp1XCQ5FACsn3rY1jdCI7Ba658wH7m9sB
AoIKU7GJc2e3hD6ogfI4vIxOAFbrFTMgZx80CJrLmMLBxroFxyx4smXEH2cBNuPv
SO68Fa/8IgGZ13T+75/juWHQH2G2/3OuB3rqM9NJs4Skm4pjzEUyukGcIbAzzAYh
bLWIrp6ZbDUelF0KulvsaY5C0BTBD2GNxlSfae7fLxtXsxtaXzJTQG8sOr5HcrVg
flK3SqaMTJzoo0lkv6JUlQDG8RmOqaeVEpSuEydxsmz3CjhrSQ9Uy3gd9AxVqfXy
qDch2cidzy73mR4PPvSraa7iMmWi3dwvFWWxQJEPf/3SB6JJJFSg+v0Ucaefvbv+
Y+bX6HN4YJbA+ALzzh7ZH4BiWOzmtb4A3wXsCK5DbzYS86IgOHg/wysNQniwMP2K
Nk4M1Zn6QjKQ7Je1fQHtk2BujWW1RCtYHVAwCIJaxcXXy8NPC3WSWsYaHAqSj5Qk
MUrlOlAWf+UxgaTDjNB7ppzqedsRDAAaaC7YuIDQGhzp4LaaOEPvES4G/sx0DVnF
kVHZMOMzTzEa/WgiR0uczdIEIq9vXa4KaSg96qY+SJFWBXE3qo2Da9v7wDxDowJQ
nq7xQ9nrLhmat/+VcT9B6C9lSXwioO6sDt9MoPawahTVsocAb5HEw1Cep0+K2iu0
G3VMTehDsqC2IxdCmi2RVxabK0/svWywQEJK0dz17GpdMzi71kCj3LEhSSNg5j8U
EpaXXSfRgnQTsSikyOYNm+fEEssAEqkzusP3P4NLHimwV9LEFaIt2f1sqmAO1RST
viETKgumAn+gUI+cv8KB36VoocWVt7FwDe0nPrhMkY5FnRYhvRMSZiq+2FCbljmx
rxVB2pWUYdLZii7SNXg0/dhxS5Jvz4WnSWv0Fm0xYy4P03Ya0NeKiV173TOVa+jj
+P9n7vrRWemIXU7CzcxUD9nCmgiB9ha2u+GXdSFtRGi8adTy+MyTbQ0MSL+thm8T
qn+xfD9McfVmrQNmOrmgqxpzx3Ru/yWDPxpMJhhOLy02LRmR0UY5PtpmWIPXc0WQ
NKGOG1n7FgegOQCwexXiSyA0Yq+Q2ejP86fd9d59V1bsF2LpNBdISYOUJLky8ikd
/k1JL3+BsMYwiqT0tE99lYGfiV/OVawyCBl5siJLe+UjnHWFk1MoNdBpLTaIw4Bl
OboxhHzdNzBzTaf4v0sUF5rBUqJNijTGKXkvrpXLyFp/cAhdc2wY1P4gOfHKMQ8J
Amr5LHbMQhzW9lmBb+e+RWHDXLdMXb0zJ4RS2mzyEV5zmgLTWcgIZHI6LsjHzdwI
P5R2KtBdQveFfkQL5CkPJEFp+9Xdmloy/tj/HbRjAV5fgfu0ZxivvwrIie+QPd4Y
X1AoDnrw5HOqJMcvo2kyYRluCpzy41nLuhD+Fl2q0QW9QrVsLcIZ76f6NNV+smnm
+JOsKdvRy7cE3OO7GowXTWSwW92Q/SBBh/m6HsXd14EVcljsVgqABGu0DI2750o0
HlV1c0CGTuxWMb1Hv6LIgHJXikCBk9EKj5dyo3KkDSwillT0zqmdzIPRaudAuuSV
XES9D1wrklsT/gUH1BW0x6yh8gwQJFi4S3922kJLFEzTHJfgEgUmiacWbfg80dgC
sbkb0SNKQX6w1y39qX1T1JQNhV5TwUhzyoyHiFPs//XjG1ZPkSujtXduBio1j+56
UkBxtr4R8bpC8n7/oRz1Vx3IhvGdpClV1P/bgeo3onATRJzz6NBa9hBauXYDXUz8
MfaNThkqRLW7c6kJ72mPogNsOLSFBG8tJzxHAxYPOo8y2sMBo40gIQul/+uECn4D
Goj2l2DeBE+0cni8JlFwjjQuhN+JUBU/soLzqtR5vtIqZBFURl/Z8b8/KtylAyFb
RrWSbfqGlyvyA5eT28eJYNjdNZTV4Sp5K+xL7uOIdWxhk/dGQwyKVaD6rXDBWVWZ
ppck6taFbG4zAgCOd68qoZ39Z5nPA9s+ZW+GD0ZCrziyER3yDDanoqtOM70xIDwf
aBFaye0wZXjx3z/x505M7xK4TE4LZ1EtJZCDJMWqPnxu481MUDWN5dnBSe1q81wX
ZnZpikrSTl6z5wxyxhPdDBeE3QLJNhPwDTGMhrxwj99sQgTkc5gJFSfda/27ZJaR
X3cfLs5EnCy+xJVI8PGv9qtUMlZ9Zmjaj3MZRfL89OMR5T80Y4tn/dJ6IgeYaZ81
hv2oFwoba+i7G/rAVWwAB/5aYcMJ9w/vJuhiyHgWU6xeeu7LsnDbN7WvsJGbIp/5
KI5ehlAUal8A0uzdfQNfs6s8Mx3KmgFnLXsoft0I1WxzKPpncc4mxcsJ++K0xYPi
DXC+Sl3WJw8msZ/MXZoIFlczQSelvrUJGSh8dkRanKqTXRtfH/hGJq+0gtmoMeii
LCFdiTsR61KtA0tk6hJ7NeOx+78oJ7FG8LZFmyU4GrWRM4ogkfv/DBoa64FPPrrZ
+jpDABE9yRMSsybIgxR0/ezUcN+Q7ZsSCeD0i1PBTK/Mye3fkQPz+4bdhb7qmqWL
t3T6mRAym1gF/XGjmECJe0h3Ty0EzrdP+8SAsXTuKyKQKSOqLHml5HRcS6NvN+J1
xiVCKdbh/ZL6cGFibpnqMjaYYdEGxYmt8TMknbOFw+hswf2Yg4Hb9F1MuIg3MwC1
GNlVijQGE65BrWmiyXjPoTeijZ5Kxk5pyPMnmG7i0g0ENyD0jfDbBj6JAp8fadlo
bUb9GMKxDer5ECwVDfz9KMwhWj2BXP+JeXUJNRyM9otGcQ2dzj+FWnZAIpF9Mmng
Sy1DfxLzfncwpKfRL6fjY09qU2USBPBGw7BIHVdTkA6vRaRzi4e/tSnmoIfBBuZX
ni6nLqOcCGO2ruiHCj3wQxa7qpIFW61SKoF0fXhAb+Lk3RvfSrv9PYJzOW3JRE4S
KjMPiDXqB9QO8GCsmJxKmPuP3Y683CYROsU2gn8H4zYFCad1ZdqwAZCqNuWSl6PQ
CRaYMl01PgbzHhDwSX4mWhkjtC7PxEg4FQR47VAqgeTydoohUwYoFmqqWj8O6f9k
hkZLKK42bPQi/je05WFifHInozSpsdV8zknUJAxtr1O56nSeGdAlF5rKeUedNXpo
Xu9yXom20GTRaQIodRV4cD5EzFiKZChAbaFTlD1uQUfDGaOhHx1US2YjIMxMkwIm
4CiBYuBZCBWsY3pUYBAXVF1aJi/5SjbySxq3lPUYudivRanvLTtiaFrDXxiPlmeD
4l6wB9vYDMkpMnU49j0en4RYsQUBdjCRoSnhegpQBmSQvnKvKN8uJuxWTI7O2T7t
znyoOuQK0XW/mc07VI71qaNRa/iN+zqU97hzJU8Md3CB9J9e4PBIaVAsvh4bsvgc
axE979tMGD3V9afV9YwbiYUfoT/aJSUO7WZu65ZpwceKCy/0mYetRo+nbS48uqRa
srxQaFlAUtFSDHd7nwj5AQcqH/PXhhEGGBGCcMhOSVnFhFOKneOv+2H5ec9zU2WP
v/1aNP02DrHQQ0EYp7zz8B/gBdWV/NUbqq7yOSYvaojnajZ/HDXNq1YS51qk2jtM
uCyjhR/+67RBaHbPOWgeUyx1d2f0IrMye4nzs3i/+OjFIVEY5u6pzAJUwkwIF/+m
L4BC8ko+giN8r43nEooKfEne35Uv3xFUDUh/fdnehHK5/X2+xbiEbGMEC6aKUkaK
Ml9gUdNrwgCeMcMxe+xCgoOmHpsde+yilwQaz8Iv2vbSWXJ4w9PDA5Dl+iDb98hJ
deBnIFuWLnNP6t0DWc45n1iTPih9UcEpiaZ3UqkGvBvSma/9jOg5DhOgce3BmnEK
u6efK5EKENvpGIMInSptTScrYMiLWYlEDjXRAd45UJV7+9j1PhCSWJ4mWN8NJISB
sKwHCLa255aYA+n3DCPWGttysFgUAZwuXJ+sfXNw4J1PCIziMEAZOcWT6l09yPeG
eFyNiX5oH4AS8EFSywKXPaa5QLhgTieEPKqfNco7SNdEplYgDlBq7Js04CTiU5Xr
sNNv0KVz77MipMDjjw5L0+0poBzdYOCKlpiTMQ5DST1lZX/8uLDjsdDDoG62khEZ
wAXCnSxlF0HxeSFKVDzBv5kOOuefDdnljRlfpvTZ4fgjS3Nj3K/TUzFw1rkmT6EW
o0Z17pwGkkBKmITwpFr1Z+hG3xp7lfhcofSlkqWPio1RJG9Dm2ulijKq6QknkaAD
g2r59oJamNGKp3x0lTB+JVN/gtIOQHQe/o/EEE8tuKkioqnjvC7qMdA4wnnCNGGw
ISYArJbCeMsbHiyR1Z+Xcm6CR4z6Do93Ifn6OUnIayLwa59C81+rSKfeIUF0LFWX
wYe1r9xFOWldNUIklDvNKhrem/RJhz9LVgRKxn6ffNAzelKcuk/iA+Tk/C3ipQNa
idXyjtrEx1/49i5FmrG8ghij55zNLRdEOftyZu0ToWnHnasWGel9++6JJjNgehkR
Du+t9tVRLou+TAI1oW0BCIeOTeRouEldND0zSZMQKQtSuZvMVNivLtPjw6ntwRXv
CPiQvbK+rq6tWbWzI+qRrpWKXAEpwT5cf72cGdphRWMmtLY+18U9YbJc2H6Qqvvo
d4gfU8wJAVq0l3H+ltE64/Mj0uqiRzQL7DRPkbgGt5rK593SCJLZUBSPOQ7gZeK9
LN/ivLVBmvrAEzA47OgMD4+4OEGUbJRGE4DVd5pUU14iluVcslp+nolJuEv42a4w
mBv7kbsYEiBY4Km1oG+r5SSgjM6Yq2csvUhtnuwshC5Js7bdlFYxmWztlUOhQg/N
MGa1sLFZnDWLB+rs11N8f9E5GFMvBs4u/NTkqqhoe5LczI1zqt/Qd25+fLc/ZNyC
6bZs2zmStgj02wTLWZuNOkFYgifEYK72+D7oKM/GkCWfWDQLBRd79aHsM+YQB06l
4ELmbDske1z8qiq15ebD4coMChoMfcNhvfSlYjzr+ZD/qbvb6pWGFcXVaDUn2/zU
jRslFygiFG1xW+5vz3OqJcsMTGO8HsGQoz/xK0nfk29NwwLetiqIrcx6GandqnXx
jYMQhh39QE9E3mKSjeiczqVAuPnqPoXlw6zqRBebYSYy8YkfqDiBXsEV/ApWv03M
R5xAD0pxyNDGMtNsv+TuE+FXnIFGWPPIh0yoFVou7ualw2hWJTB8Az9DaKAeP+JN
aYiOo5FueKujtZykSanmmR58o0bHfvkN72F90VdMBPaVa2tMkTs+VwLHmEMjAX1+
1UIfZnHXoo/u0CuS4kS8V5vHEgY7nCaHaG5FBMiff2THGak3TwvECpLBd7gEhaGh
9ZQ8KosrSbcXFM6lGtMk10FKGK+jpAhLWNeRb2GMKHK27Va0GHhCXKAbXO7kzN1Q
nCkks8wZqSM1rtW4VCNFjArZE5R9iI7WNrJuKIuK5y2+g/4yuqnm8qvmMQ5KQ4E5
2M5LuFpM0Nl/A5hDbAhcMfdzwxVfbxT4kXFtlo2B2qOkv9z+oVMHIglsm35CVWk7
IbT9fUx/a952bFl2pZpqJFuG9/FrJZ2/rvVwwn08FUc5C/5hm+RYrsql8+J6Pj/4
wex7mcQ5yqpkBFELc8mN8IrNE2qbNBWn68iqga3Rboo6UlCdSiVA4Da6B0Ddp1jZ
0gUcLev/a6OSi8shxSRia8yO/KH5xJE2H/OLdwmVI9sO6s89iY/20Sh1TLsdCdZf
yJT4RWIuk/6YI7hmnDULfTdbvoxU9NXoYmg5dh9A1VGzKg1cPsE9/LCQx0IU6xL8
JV51PbWbG+fI0aJr9FrA7RZt2GVg6qwVG1nEI99FHAgn0uedy+A8PpWRgi36jZOe
ZhRHP5imxEykXZELjgF/dYFtLtOpWofrHzY72pSZqHuMhkApw3itz06JlMLJt3ci
8JAtvnM5iC6KuSQXe7qWl3N7MXL4xPGbSoEgYXsgBgWLGDLU126Lm5mtWKF6veYS
6KkTHQA72h1bL2PsIPJjC50iqeHDSWzl510Mmq3csdEhSbPHk46HsljKOr5PgxrN
HpAJfQWrNcRhyM+JJ8cY8hgVVEme0UEqTRlFL7SwO/k05afC9eC0tmxgH41BUl7A
Apb09mybQILX1E2942HNwaaIUrGVAjv821ZHi+wIRCBXFpBC+I4ti3CwZn8wkBpF
LHD/BLyH3kCAmexg4+xSGpQaDJZxwHqlPaloaJDNgF5864mDdyV9lrvRSMdyNcmF
ImHf+JGOz7uRnoSdQHa/9BlBaBAI7o2ZoaA1km5mLD2ZCZw77KNX69hHDS6I4gDq
maRm8os30+VOtqHovke1O4ss2lYqSG1WTNg1LXz2im3/8uCeUZ1pcxyIEqwTlrVG
s1AP1+388tcowne8Tb8FMeR7KLARzWmFui9nsJuiPXRA/eTIcyVY294WNYNAShLy
3OKWqjXe7mrb/PpxZbd42YYur4jISzmP/ocT2gU++u9DOsGcoicJ0XhV1TAF4q09
Pc+0TIRzUJqkRlcUbEUZTLXKHBkFRVOPdCbiThem2NKGGXa4E9+jLtztLUHsg22m
UGyqDN3EvgOe1d9+iQOoKxrsQ2ytZe0NMaCAghqqHSJmRujm0st1nS9oJjk7UHYE
QL0dyd1UUFjnNMs8aBFHxpRq9nSKh3Hw6fhBVKwmn7U4BCTBYIDKaxCbuQ1+EmFV
JheisPDIuvmWOG0+6HNTOUT6SMSlEZNRwDYa630qyZNvlxA4HKsys6Iuvk6XRWoa
+VZ6SD3uN0brs6woYr5OU6AauVoZv64xQEz5otp08NB2HmIbNoPQpQVDDfWkUS5e
ZvXKrHLbyBQJflOPubI/VrbKIftyHKq1mkr4ZOBD2X4W0kuLp8F+daRZwMiIM6zl
LwP49+ukYef66isxm6GHW1Ew3JiwdkKInUnTHyOlwgOrDVE9ggrXdUR3zl6dxP+L
13z7zBkZH4xehWZDDEphN4weGMpso1EHeavqwg1AO27DoBE3QUVcal/S8xQzsfBM
W8lOlIotJJv/s0YBWNgvwgfKIPtOyQBTQUWp0qe/Qm0WhkLrM/8orbutEgw049ac
KFu7dclA0U6y6zdWgByV+gj98rqegDoYZsKuPYO7jpCNqgEFzKEV1GZFUBSg0Iq4
i2/kbPbjzvLhXyHE43b9HEJ2BItVu/XhJtcmWQUn6Bz1qNdutdLuMbPTqYl4u1qm
wBJeboUF6FHcJoz6GS/lSOKSyvnDZKMpYoyL4pKzWoiASY2UcEKJ1cwkWrsnLazJ
dEH6TQDfMX1mQ5YpwN82OgKOfKL0U4obeTnGO9fDu+m00Op9bEkzFLLyuINnJiW/
czVfvj+yWB67BOBS/27sH9Hk6dqwxlSKstWcLCAcF16X5Y68zf6fJPvzLS4mtWdO
0lBkeLza1Bnqo+YhDw0bGdXawgxWJ1FVPc//D1Qg54G6MIw/dLsA1ZiAhW2W3z0m
ibAwDjV2rQREfyaP4Uuylq8HFwVhCKYrB6lXjVtu+TAwtmcx2lmjy1fkpN7xNmxz
KjiACr4p/c5T1DiJJWpUkmhoaRReklAmLip+o7SLx/kWsLCBT8pGmiKVFmZXceiX
bLrEnbhbKDnfnvrOZxtnZtvFg+Go5DYN/XmDEICefdVVNHj8Lzxs6nX4uAcYM6/P
zl49evWseQSkQ06i+/ZEC2VW0yUUlVGQNgCy0DaSBUeuN79WYvda0W/Uvm+IFq9u
40prmQNyLTc9XV+ZS3uEsRgf+cSPooNTfBaRHngcg1yoLfMamKZpKW8mcOFkziMk
1IYRIEHwcJtIMQ39hGSHMYxrZSnGHqHUEFO47NMUeTueWvooth2amnBSEBlf67pE
qyLD11EpEQMlCoFoWtRRbPLXX/ksLhfe+iWcxWC1cytoqfdhGBj9AK+ZjkODERVC
T7V0BDssgQZAQH6jbmfQw99qBU47m4UzUscuJXS4plP0hb4jkXbhSbGhARfQaU1N
0BAe6HuEBUvWByJG49JI3ItY3bbGapRU9XtZnJFCVSmUwsM1DfVJf4xHVK1yUJOY
9uiEuw0yawPp2PEY0hpoazK9B8O8D29qguFA5uyctBpEjevVFkGp/82BkTZ00rPK
r5G0KLLsGoHBgS+kD1bAEPhbevZwosQ12shUCz2SuIq81ia+yEW/UVa5h2hC4jPv
PRs7fnNQ5G9hVL5E+QOIyoZE2t8tk5+aAC/Q3T5ERshf1N/BV0AZqw1UXMiFywjU
ORxK0PFWT+YSAGIqmQXladXXy+4TH8dAvbNjmqitS7kYk/7jvio2uBEBzz6Rq0P7
0Fef7TBjzSAdDDp3zr55pHILe0q2A9uX7Lo4vwDMqrsaUdwJ4ki/sn3xvw32qS6y
LRqyfxX38opiPvoBQ+65+EA/yX5DFPQcWdwOXxMvPfhaGZV9+ZcwjcNYPXAtt+sa
64gN4dVm8vbCQCWsYeAN7h8BnXnpP0Uqa+wnoKmnkDC86r5b32Zk2A94W0/MIroO
D8auIZtz1viu8cZmyHCXLH60Wwh0Mkr/SPPZ5ByU1seMlhLExV4oSSMnFg99UkNM
81lClncg60bITpzCqupqCNzXN2Oy6TJJdORMbezNTFtK7fEkzl/nKuJYfLEYzoXB
Co4bofEt6LDEyhWUqozjKGSjdOKREvSRp2ygS+1+EqfFrs9Pp8/WxmDH7XZ8Xr1l
UvmD/1JrN8tO38z40nNsLvwdbeNxXNVo4kLxDt4NL/4SXk4Ml4TYlOL7Pf/IagZx
Q/xy9PDFBrvIQTWAbH/3eKCkwHFbOHg/cb2lUkC9FK6NpWzL9nzlUA//MnP/BsD0
vRW72EHm9Vs9F+OO82tKeSknTXFKmnibCC5Y/1zpxH4oQT4eHI0TETf9A5ey8lW6
T+FcDCysbFDhlAUtcPUySUr8dHED3US0MOsvnDGKy+WlKTM+ajqoqzO3omHRuuOz
IR7s9NJwED+Xc4OfNokkKgWNyWFwLsuCJCz8MJO8y6qDW6g2BFZNyZBtZyKq/t7G
DCuEvBBBIHQnJdSdEhyDdrfCg/2j3O7Ebrq4aVEAttTPmkbz57bZww6ydxP3rz70
V3fw34ts42U63KCiCMe+Mv5VmW4uHntUjGc0jrydcgsAvuxqUpYbuOHOwZGfOTr5
TqGqTpuFzBsy42zU+JrbTmengQVApSpynaWfGf8/4RtTjz4pc5KRjYovMDXeF7Pg
HzugyxIqSirFaie1lRuufT9mplC5u+LKDYKzpyrcjdWa34WuORpDm695Ap0umReC
BP7DPG+lEDskO1u0NPs9thXBnWH7WrZikeNUMVUOFiEM1pgBNfCmsHJw45LDwSya
jdNLxruFKS2d+TfaJNpuaurQzLX39eFWD0VZS2ZmmAV5m+L+R9OYZ8SaFFepab/D
K4m6m5F4jQIBrqVqzXJQ4NpIcoYXRjKx6UbO0sLVifmSsJ4aGwiYP/Pmz3Ts9T3J
uAUvCc6ZFGIa88NsnoONZ+uafgIbjzWIzXNcblR8sJSzu73Ce3f6Hqfli8vJVg+g
qjrPfoaO/CAXb3AcFDVAThlNxth+Z8tso7rzQH8FyoV7DguIq3y/Zt3M9SWhvscd
WJdMwp7RpgpK7sZMOuCabZxMZEoLJmQJwWqaJWpjOrR+BqTEE1qnIsg+k8bsMDME
iReDZ+qLuET7w+Glyf3SI7qpwvWxcyT8iNthBqOIWFgaE9naM2A3FrD8EBtsmmmp
e8es2BIiko2Bu+KWHyFXW+OkdCuNIn9Fg0hSuZYGv/DTs9bccXbbvVbrBrSFvPIP
pTh9wcYWxL3qTyw90AK4vOCtPjqdtaGV5urAWmv1WDy++N5V8UlmIBXxt18OFb0X
7rWlXlSF9XxkRIu7V43s4t8pYof2JlWJeb30+wo4GJbdEMCWVyPTHGjvYvewHox/
26KzWUcvXbLQbZNmfNX2vney9a+7ouJvx0XJFv36FN+HPhX30cJGzNsinPHar4U6
is+UNAb6oRvqD25CnFTlxScpxlCyT54VMcTazYgPS3zPe/pG5go8hk02VEGUdy3o
DnEhAbVLK49Q7fpWxAZKjmZoZUhL2LCHfTaZ7IG+JVkVOBAf1jvZ3WU4pBvLe8Em
4fH8U4s5mLVd/XbTtVzDP3QT4G9CRzdpCl6spcg3+KTuhmLF/Mb5R6UzYGa49Rgr
YQrL4W+VZ6gMIJGx7ARAe5YCEhTVr+EPnE8h3kI2ieqTxQouu58syLCIO7HxjuLB
a666dSv6VfpMKhh1i1riLS186V4h2tdC7EpNW7kgC8VSNCMbEkfCc0IYx70c68Sf
97wFvlqAL6VTL+8eWFM3eZqNoOgyUNh/7GOsChgZbdfe0Vv//lDEY5pJINm074ej
SdHtzyql/542nr1Wk+8zscGMeXr7pU4ttdDueCV2kjWCnNcECt0sEMCjRBA0bthX
83mxnqaLLB7Kjc/VokJAm7flzXuRskDqu5ODhdWrF86DJDR0S2zjSma3qnTP8l/k
3lI+UmIfkoGT65b5pMbX3yuFIYSDehj/1ON0MJ/IVBiMZXdbXwQ1MevktvOQ/y2j
3kk2klgj+Y2Csg0NAY4lauk0zD57xwoXlNOyamtAAahHru3yRsMow34ArNgmAjtj
qQ7FPwN4urz2GLWRmvPzgSvVq9DGIo25EYAA4ti7mkhjILd+xAiII87GWQVDoeIp
I7yLIfRhp6WCmnbIAoOPeGsxsBLT775dSTG6cC7YBQjYmCTHZq7BwKgsFHsvjRLZ
Q7uoY9G1/DQDfX1cItXI5IqCzZb+Rljvkf/DeCQeLUIyA9shcIV9p2lDcMQYZclt
A1nz222KVGg1riT783js+ks2meYPWGtsPOlGQfSEG2OW25KxF0ns4FFBpSs1paPQ
YkTddX2zh6qrBzSqw2T1/8Aft6JM/dH08SwIYSvJclYkalH3MX78bli1NBy/O6aj
RVAsvVPKZdWWOlUEQfUfY6lBQY28S9Po5BMtqO/gxLvLGKEhM2rHClmGeprpW92G
+KPWwgxV4lSO5sy9B9ID0YyRxMgWvJkqH9hXD0vMZ3OYCewn8Ne9QVQZkkF0DGIH
S5pWXW6ktJqzUKjtYAg2S5RiblWcCeiKWTFUZ6Gsdq/KqdPqTTk1xvA5MvHbfO9m
IOEKUhEq6inlyZ6mC1nz86SWBpqiZkvk9+tDkwB0cua59duzA+gdj5FG9vEzXQr3
R/ZtliqSfumK2DomLTk6LB52fqblZfs1yQDaNaLLNC26eCv1gSciYPcD9h19ultl
sX6PJi3cQ1Vo9YdsT0bvFNfr/YzTKQ+Lpv2x5nZ5ZfgBOY1n1EwoUIFmf9IIWf/F
17bNNz9oCMrcJlxxaFV+8rJHby/A+3FRbMZ6U2rCnswCn5Yy4Ohyv+izK/usrA9v
JkdhVG652HsNR/iStLpGh22AVR+QgiZXHvDMNF6FlfKT7W4P7oLnQNZLDoxBC947
3nInasVZPPyOis1BDGn0GDly4jMw/XFTtHbh7dLy+YJgPFWtkQmbhTytnYgHomRn
Cm6PZnipNR/W9mA7KEvreJ0bzyFi8XZ40Z+HXy1/Dt52q7gaG8AhaMNRsoejjhiI
yYiMqiRQRzKm0bqPedC1id7drv0xcF+DfMwId0F/o9Lx9vrGsgdZbRnvhPrA+e6a
afj/26siIaxXuatWDmgMksx+BkD5jyYVk9d+qkPczZ+q26RsWYJK0QPfWw/off8U
/YN36vmL4km+Ri49uKcNGLSMin0ec25hWVLrCG4URwtNpVTEY+eFbVBC8vxG0bxL
nFQNIGYOnAMWjOMuNnEud/vElsX+HUWeelvzGcB/0Z1Cn8LQ6y4wBSp6ZwzXHPRC
UWjJgqG2Tej4QubvjMp/j3N/NNjrlUt+YsgoF6c7gwVKRTnWmKbaX5kCakOU/URq
IuTFcsICQ0LHb3tnYMfVfXJNJrPIDF01kHgKs9Fc4Wcl1pOViPOYloNjUEIaybQi
Gw26fefyltyzOZQdFI4G4esQxwthaOgaPG4E7ll3f3gstP5gvgk09qZm4CUhzMf+
4Aw43LVXCfhBGW5pcfaaEK+lphQmfckdDZ/F24xuJuX+S9W6tdbtmfXX1gZPXdyB
fvB9YkzVbpRS4JH+3jxLZQafJPxvtWAlEUPpyIenYO/JPYYsmd+9uH4iSLN+AGsv
6HqD+4PS5ecb7MjWFT6eaChcZ5SpDvGjaIlC9/obZSMnQavsJ2axk236MfqS14/m
3qD2asSGtpBas8MdiQ/VjV7AZORGDC9Jku5XW0Wiu7cL9qsbMyvV9NaHDnc1frE8
H1SxfiH5v4pEnwhlg7OpWd1USGhIZa8S2ylnJk6QRjbR+roV3dBsRXAfnrM4OfB8
F1CPSVS/xmBlygle/Cs8rriE9XvvL+dia/KwcCSL04UbQUswrMFCAm6MprTQFeIT
8DW4uZmVJlIibhtZhFEP0TehvAnZFWcylisInsiGmZQSqe0uQxtoByi4YO8LApl3
g5PwkKnFf1IXDFH+mYHdyybZ4tfQ8IdXuMY9Kp4jjDRtMQsJL3p3ba81N/5VF8iq
EmEPhYGWTSYrDHhHagjn817/ZHHYGL5WMxAoTL4rRztnvngc+5nGrsBUUt4ktLKK
T1xIxxNTUjXURgCEbagsr49Pf3wW/fH1A5d5Nx9rhIUfonsvA4rcDFiQmOe3tmV2
R69JCSMk/ZIxNYeyV++cZGIppUhpQmybjbl4X+edPQODcOFw8YG1/SCdtE3Dcw17
LqdvOs6Hp9UHoL5EpTLXOBfXwJLv2HcuaYXjV1Axxel5iXLFFhehQdAcR3pOcc8k
bxY4L7rQX05k2nI7kePWsTNyRbkYxlDeILnrOG6H9zybHvt/QOIFaPP7QQsJwqnk
/gQY/20MDmB2Rf3VN5uoKS4f/gWvW2ZJmOO934/UZ5GoRkgemLJUbPvalDo1dUdn
4f2yo3jaNnGFXePocLuEd47joaI+ASrdXCDeVx45ugXi+WDNj4q1gSj0axESf/GK
Z/6kuB9FSJpKTtkWzeKybbfrdUrKEVma7bUUSBEC35pZKwOyo5/FZ1XC7OeNcwZO
zJ9e1LvC3itwPj90FoUOLQfCh6AIM/2LMg2e89F/ITMjnlsIR8jpmzt21K7S0Nad
0CZyDPTGY27uB2Oq8N0/+C/auAWDyLspHkyPt47n77yBNTn02bZSS50Ja1aCjhn1
2f5gjPj8tXKTO8e7/v+3BGju+R6scBeing01kwCOiiOoWLGMciKi4Gp127hX/nTt
yy/pJ4/8MKKlTsT2jd5SldSEkjydZ0Ob5OkBKg6flfnvOLmyXEohJYxM9Hyf/A2A
bWa/Rzv/pYK5OXeltKwARRMhcPGfs1hZifV93RNK9hOY9N6nYKTVhXbD+Ng+YQt7
6hMLJY6ePMk1lK+AOSmNs1GnZHvYJTFCW/sHDbZRAkFTy7yUCQVI35DqogNORjRy
TqsrNhEe+d6Fh3ajNavJS1GGkvTru7CPNEs6mE7lIRlSiK6V7zQTWoATl+fjLzFr
a25q4Az8QW6WAqEHoCXUzA8s/eQ0x9IinbErov2mObGz+BamNVtCSisU/DbDoshs
teKup04jgeT/rUaC5GLCxVzKf7VmRLd4Bily3KMtz7NihS/SZQh9d0ZWjekZxK3b
WcnqmtPAo76HUEGIQBSS3WGGCtr+kfL2JPJe0xV6AY7oi/UQ5uYL3E+MTkmzYS3l
ZdRjR56M/ICDtSjYMmDeO57nghnO7NHELCa4V/+ALiE/4ZWESF6TA+SHPoYezWoe
e0FtWr1q5PXF30hCnm4ptWaRsxeSpWl37ybgEp2vRf2ed7a5wiKK8gAIpoN0BO+5
BpnNGX2Z6tB6JDdaR6gy8DsPVUI0oULjydKtj6wftnKSvadN33clONwIh9oOVi3+
unb+cCZVKa/UbCG/Rsp+opo218sV5AMv9bdPlLxA+HCGfKvX73h1fiu7p2WB+AbM
8v8b3hgYCLtffnDdJvw8qGc5df+NVXKDv+r9E6HqvFsfxxIy5x5NtgEgcW3bkOr5
lvqDOMXGazI7hYQVMk/ReUJouaJV0GJQrzhhg5sdjPCgZ5ybYp4XvouiKYKr0jWS
SCRD1x0SFtlNlUgD8OWhfNXiI7UTO4/xyiK2+qzT+eZRQPDFYPK3sdL2DMNXNgRD
Buh0yhXAJy1JZ/ldsEu2KweXuknxAojJ4CpqNN183H/m5yihvLbOV3lILuUaYHxh
6uIfLiadDsFffO7Vc3rWtGDYqm7I7IGXAaFcx3RB00QEdKoXCAdbtEoKsHzAp+M8
nvUX8bf/lu7BjFLrYvrK5Gt1nNYXSISi0PZxtRpmjqG0lwNUImFgoW+w2m0+0Q3Y
bA4sPF3DenrTyf7IBzEZHes4p+gHgbPivkhs4A5n2+HUcrCF3dmRZT2Nhe54UYkz
pwG0Rbppg2U1cKeTEy+927x7GPM1CRbqaXCOU1cQEcT7ztb5xt49Pusk4P6BlVlg
a/bqo8uVz9OI3J/ZmRLlvhaV0Lj/eRTTU0EIDHCI77zxaMDjTpEaZk9MqG3IPNX7
QtM+kp3M+DC8/7B2rXl8nnUp6AiKtOiiGoTkFlX3mLEPBwIFGkfoJ7YgqJxyH8O4
qeDhb3jeK4mQvFSn+w6qH6lJxCtrqCpnLVQQT8bDpGVfRpCtZkv/MrUn1zje62mY
hPs8qjYq7AVg9aW3jTETMAPJ9oC0pj6ChBHnZTr4BSG657RWmJ+SxX6krtR8Z2Wt
O6KjyigO6dndY9UtzVIJNgDaY/rwbNM+IHyAYPw4dbulzxdBfOM1MwR6N9+nfkPM
JWocE0qMAwo1PCZig7MkQDbB4aqIydNXj6J0V9YY4IUmo7Hm1dJDo1z3k2IiNrcO
yY9/ia4teETKMwg5xf7JPqbXDAb7heXLP/pn9Qvs32Hejxux64jioz299/igMFeE
6aY+KUETOVRYLr7zAF6l1Krxy243zg/507rLmykjj9orQc032+QyX/yeDM6n+Qi4
uuv1h77C4eLpJqMrV/MybWr3b38iK/uTbcr2KYjIX3uQxe1Ey4a9OG7fySjbzBcE
5eOyDKI/mMEljLqO8NnwKjCGYf/pPqBwKSK9D7B5dsi8ldche/JGVIaZ7nUfH85g
JJOUH4+uNhU6ncCmt+HDSms0BxRy3lIxItiXriVlv0no96wXTUQMr0Rn8NKkNSZP
TEpt291DaTxMHkRRAEa+amWMgmhhpkvXA/C9DiGrZrea+OA6s9BZ2pBc7luGwHE5
XiMvZedyo7HRm2PHCkTzsEgBQJm0cMJvaNZMc0EuTCsBC8PUy7JhfrGW/Dwer3Rt
OsMLu/1eCZvf9rkRDyjTM7ZOZxtO3Q/UEnApMwNbSpPCXIMSHBu1AnbJ504klNau
7hUD09dGwM2BVVOjUbB67i+y5RfYOtuVhHOTOUfsxv96a23lBoGUwoxmPmyJIWGZ
CBzeaAChKqr2TmJF5KTkaPmNxNqzpcL1nPCLQ1xfxDBCsTcNPnXXSQ67iTGi4a9M
elNWoIRcUGlWYqjgoPk6nFSYDQT7wpeizBtonE3C9sCJhbDznoCLj3MGdC1q2d+l
aQkdQNd1dMXq5gfxU6wySSsrSPPh8Vi82AGULJ5+tcbmThJtkzIKRBFvVo8BR9DF
R8hSKK5dKwd9y5/4Icnk6OVFKRTviqnrYRQdFFO1XiWNHhUvP0AETFb7hyhk0F2E
1epIhIF+Tjnkk1e6yGSubI3knCQwIXw2d1hAAvSP5qXqVNoH0o63J7R/epC5wvff
tkdIQwYpSjYUY0iF4Dq4LN5mIkQNUC7ldofIaoHD1vm8SLDw0Ld/f9DDAvA/mGrU
jARZKNKy5b8+0jVsDhpr/k/IaMX08bHYnXiDpD+ERaWabR8PKE8dc6cAQnu1I34t
XEIhom7Vuk2fOErc/nlEcajHoUGCvJFNgLyqnqCwKScay/G1Tn0+axP/UVs6o0DJ
FPh28pJXXW9V9Z5W7OkCouxevvJCOg3Q9+5v7NNkaqPV5m9XHFKLmzbapHkx3Cnn
23SibnE2v3W21yIuvBuyUCRKiPJTEka6TDdzj2c3iR/izPKHxRczDTW9aRyLFq9a
EjBTqaH3DXqY/GvZBdIkM48NGRDeKkwU/Yn0h78U+VkeYCyuJKVm81Zor/aOFOoJ
5eFuAL8cjd1HMbMHzscHBd7kqh2Yo3mX0SqSZUstslEcHApr27go384fFtjDyMl4
8f94VgytuID1Xyw0RlmOkuKQDynZPhwbfm9yI6hpvTTATYXsaZRFHuogg/S1m396
8KA9usa7wW56mXw722tV7MeXch8bUD9T6ONOYrjYPvWpa6/9qvRSa5ATs60eOD7r
XMN6fEi71zzxNNdjeJIHqpiV3iwq1eIKGW8zK2Wey4YXZ2s7HVNlLoktjQWNmmKw
RdZGaFblrwgmm70uazbPW6tZv1hNJj67L1pWxlyHfPlYT6WjaXFT/QYw7UWuNfTM
gyv2q9WfCKpQnbvXR6SpIDByCwmEvQwQ1eAh0JRCRu4wLAP2/r+mRJmdVtKC8Aje
Odu77vqqDWe26kpbPIF/gSNQ1p0ePgRzmVlkIaewMhN0lFOGOtXid/c3LdDpmJ39
rfBDYUCLzLwsucwjZJqN2TL/RuI1tAqdOVtECmFH+5e/oM20dbCqBcg7y96eXOoT
jGRD4iv8qlGZMzTT7AZzTFBM1FiX8tJs580KdM10GuTPCfSubr7jL5PxQznQDwwc
IyOFSBpyX/yTaxKqyb0U0a0sCaAEZYr4J/u8F8nyipKx1YW7GTCx8TY/aBOaf+bK
qzc9+AuWzzr8SxTtOyrxPEiHT7Fho0GkSQXnK9wL/8Bj03TrvSWFyp8ikGrCgIHL
Zp1kb6OMCf6uvVW7ITFnszPviA2GtDgEmu1j+pz7MDXTdrt5W4phNQb7LtheSh9K
huHQspGAoTuHWuPkVhgd97Uf21pvJx1/R2AdRwZyJhjXO90o6P+oe625dI3ZrUL0
73pIXi/ugFSXPtoV5WLYQIQXlJ4LT4EuE6lkigcfQR/keocOch1spaweoNZaDEWA
AQPhXocK0/D3VHRf30nmOlavEuB40mWkzNwnq7m3vNvqMRdHxlJVZwqdRIKYlk1P
1VkOZuOy8bPtYlJXN2Akdr2GxovSjfNeZ15o3cDsarQHXt+2WjfhWBH9Fe0ofNaF
6/H2JCYyrC4ftm01tVusjTGguh6A9z2StjxHF+2s5ifo9Alqqo8+FLgOjEIajFLG
9wGKw+SntqsiOjnt5skWH5tCD+Vq66Qqp5eGqbOKZBwU7wHBUwrNCmWi+EH+agHB
dNmfU3a0VkzyhuX09tRIIL7GO9pVIA6YS6v/sljEie8AQlV17RHQmcNIcweiKQFb
TUIlFqG1Ug4GeOBjtr2EfdjYnZnKwn23jGYMIUb57YsKD52SQ2kdPbnqge1vxIXz
mHGXJkU+0aThuFAJZ9y8U/ejyvOTzhCHDvvPrJvXHYqz4LeHjxL5xgULBo9LwIJm
qRjZy/ANzldmZ8O1YnyBVE2ngvdAc0yx79oSglc+mTjH3vRzKOjjhtBFiKlHAt5M
qtvIhaWFOZK1pX9K4lC4FSo++ZzjqInkTgpspIrasGjzHVdmfQZoFdPilxw1G4wH
Fq7wgF94WExMmusCL4BQdXueFUl0iRC3bzpf1nt6297u1U99J4A7EA5vV8W1ivCT
3XKJYyuAcd/lp59/4jVv+OLW3ZOFjEhMMTdUfBsRs/4tgm/SMRcJc6DpCtWviZcW
lnArb66YK49jxmAK0irlaYMUyrXpIZ6Wyausc2lQj+WOdkiu62bYb/MjBnj89eqF
mR9YkAZUuhcOvGlet1sa8j+ZE3GQR+rAU1g7WILdck4wjBiG1GYgslhzQ0nY7A/r
ndy8HPlqT1bp8zqZgCP7Cre+K4mtL/eZ8qKiZR4UqwuMG52xt/JwMfMajuOmhRmD
s9ElpbwYL15j8/2Tgd/2NTDMsRlQJyFmkVM+ecfCkDSWcUEBvq/ysh6DSEf7p5D6
cwH5zhiNMkp5//ws3bHg6fTIlriS8gWv1tWzZxN6oNX/GsUgGloeSqOMI9LYrItG
aqNf2hEF2DO7RBBLXyT6NvD8T3eiFUaXVxd6iuXHngfW7uslNzlydURnMj54LH0X
jMcZB2aSr829UctkApyJ49kYyHjyrcDImrE+uIG99TPlA2o14el40uRa06rQ5A8/
gLU4e2m8cVicBHdP010jqYeCaN/9/LPDnYmxJoColTTBUX+3XMDLtGa6QMMp3a7J
3BOUFF3KWS4FfdqaJxIpH069/9TKLHwB+dlbmVrSG0y+1c5tANNxaTJf1S4EswBJ
cewzl2SMDXUNBa0tzL6yNZbzpfTjdF3pD19NOXSgcjLqG+SuHUffXiQrfnRPXKEH
gXmzyVh4M7riEI8azJglNKX2M3CGOb+six4FzWpqiO18/Q6igINWprZSZHzsf0KC
eGM1FEfbGY1j1VXTYfWoKQ9KJDPj/eSa8XwbpgGFD+lZq8baiOd++bk7ZoUnYqzG
uAQC7vNI6D7htWgvhVsBvQZZpb/JLMrymM4mZ5D59iq4Z+YP+xgq5fcpTW3NHUs3
H3PXG1umpWbNlnBNPOps9gk/hA46MJjUWPmZz3wDulyRqRpzGNtoonAMltopTr9n
b4ketiRu/7UBYBGAZIfPJp8hu8RE4/SHA7bNGvlTge8xXvcGlMwUQos/DdBSl3HF
LrKLMV3Bk2qYT1afDwGzXzbnjAyDBOI1bTTMqHO9FbvsnqsH7qQo7X06xtNXA3ui
3mtxAPosNj+qvdPDuSccADUkE32Jb2So8gkD4AfCnofhe62sYTY0SalQXFqupT4S
86a4J+vrMEhzFz9oCmTD+GAJp8hUN+z6HTiWfR7qD93izE4UZIlhGVXA7giMestB
Z8xcAKszn9OFg1UHsqHwTv4vvRfOAgzLcfaCjn54Dy9dtNvqjxCBnCXpmh74z9O/
as+PlSisaw5fwW0IyMCJNppwJztoVJxiZerUAQAPV1RAvG1t1Xekd+1FAzhMZO1N
esZKX6I65Q1M+EffYVL0sQtyiU/DLXDJaHvAZzzeOkUpGTujPhB87LDnMtWSJfHt
icJNQEk1bpnko8AOYbPwNXYCeDGhjr16IRq6j+dcXpxpAupnhX6z/j8vKwjP864C
NRQ1SBgMuLQJ2dClDJkUsc07C8OlZCo55GwmEomFUnRXeqmig67BJA3fIMquzTZK
B1nyXrhL79S+9+NpX3NvDnJ7ZSl7NzT00XcHE/akwE0jqsRE4MqiUeY525cD0apB
cvPoAdO/RICwH2cURcNZqGmyKJyx6LyZ/tdBYSvp3ZhBOrDsUj/sDzuJtsigSFw9
xAtO5psaTYDoQZR2vmMRSX0Z64SZUZGhARWFgrZSoPUMLwSZLC0sgPJvyeiKLIsj
Dcw7Kz7YL4ifZAM7YPgWO/nNTMqwcPrQrqBH8QqL63fNlp43gK4Njw+FRTkINh5J
rBi+GuTmyJhMt8aH8wDU69q+8KeVDLjsPMsOSG/KbD/ol78Ke3gftv90HUQzRxuE
eUHRopQNJ9kzy91fsUwHfC0G+Noe9MgvLpmzwKJLB/S4hCTtrenZifBf5HLbWt6O
lqBOc1GJJcudr2peYx5uMtdR9vpPhPgWhvvDzKoTVAVVoca0Z4CW9bhVy19NCz3W
BLZqfo8b3ShsXaRjUZIorPKrX51nritXdpMEDUtnaG3PlINOMoSZgbRqYXEHXO8J
ZvU4uCn0AbaQu9EPlsoMenWnaPs+0lpW7NHLju7qyMPNbLeKe9qxIG9xPh8Q0gaP
GsM7dgH9Xl/dZAEWrF/Zqku+4KuXrl/2KIw2L+Q2GXAmxZIZUhnxMLWQ3f3KGTJl
ptVFOOpwIJDH4XKPQyyn6MCHP4hzjM8gRJtphZG124USBmzaZrwZnUuRsTZeZBeV
FS6LOoZTqtS0W5f0L6mrUXETVVEC25NJi1EHGpo9jrriXljrdjZEP37l9Rck+r3v
6yfBPvff4oT5iYHd/bAKi+dOJlxxILc8yQ6alPfWgGpQeVoMYrup6eGbhCxTadGL
FQYFROcRufR4bje5bx8U98u8KRjLyRDokWvJQhhf2g15fmLmRbhRYshSY0FX6weX
iUt3y5Z+UPxiMTKIU3QdqiDEL7j1snXs+dqTgVQw0kWYOTOcFxcaOHaO7JRuXek1
7cwM1L/4evqd/2cPko8xo8DrEr4hvycap1irFGw88jxYV998XClVm5zcRVFj0Xgh
lztqhbAfaLZRdAxSd3KGNiOegYZslynMEVkNSL1gA685i7BVXvqiKr+e1iO1trMJ
VeWyP0N9I0itxBREqfAaRhRmq7b48YlmaKkTj8WmZjilmubrhZUrNw1j6ZU7FXBv
0HKSJdLv68hwOwFtfHwS5Q3A5P3SvjAs343evbYipIpYKjLGgCHgsOrDo2rzmryb
Wx6bL6SBJEY7Myjioe5NR2BBckOZaI2rTpWLVEJo1TcK5m/32hTUf6AOyz/Tfq2X
tofv0zDqL4/YDMrnAaMHi5iOSVclNI+LlQNqHYw1pg4t/LSyomoGLikrXxGRUsOE
IPMmTGDBLLInZzEYv23O6p70vXRi66V2wX1tODeZFwN7iSqtVZMfqeS4YIHTXRwx
qt63c2iEoWFl6tLRPcirjNyMJFHQjrrA1rWZH4LsSImcCRXpS1koqL0E6O40YXrp
cG9syx8T/gHmGGlqo8JIrYUWqjOjfaluelPbEALO6YiG53Ihfv+Dh3MuNDOSAtJ7
D+ttAhnzzgZIlurxuXrvmg0IZUP4oRi3CctHNCIHkH0LQpYdein182b2k7iTsA5Y
gt//oV6DZzkIvNc+weA8ZwM070u0eV6seHmJCSm+iQzBJ+5eNxSM/M6aGAaDGCxB
w43bEz/1MOn73B+KQLEm15H8IosvHJlBcWaS/paq/kTh8KkX/Vs05hW6tlv3DhMD
b5rLtpOBMEkxQW1mFUdlUJWlTCoZ4u4/n53NlhEpOWT2Cmjgy36o49HGC7OUP5Ed
XRkI3zW2T5Qect+s1SE3uhPjb4OBb17ZH0exPiBPXLBo7hhoM07GH3m3xt5p8ccw
EU06XedsVhiwC+VYMYRSerzffGW4xxpTKhegEY2w8LhKQyR6FTEj9T91DctmVEKw
hPezqQ79wAkQwdLCOhVggehakN9wgtkpvDBoJ4JkXdPt6yE8y96uki4rizubPCXu
LYewniuB0vh44BbE3DHSETQbqRIEZKAZSAya8M+6tgFWIgpIqbAAweKVtWKPhOSu
7lqGHS7sKiDJCXNNec+u7K4KA5c47qcZGFrbmXWlvzC/Fs4JtGApwg/KEnl23MMf
M6y5kXFV2gqheP6nAJkny/j9ltuUNBMcPZfQ6GWFYSgBDmbiOqxXekWeqJSEiLnE
Yu+YxRDQWPLF+W/c9gJ5JdJo0HyYIXPj9PQhbcN+cOf72HvKHegBEy97bnvgct3K
/xNMlEp813qmCp783UoXUsGKR3KtAlzg2yU0nuBLWF/E1ewAl+87mjtq6sniNpPt
4OR2sBphcZt36Fnhi/LQaOUJCPsrnIGDedtF5BVDlUYKh0Sv/6yb1W3NhdpuI3dJ
mLbTXI/U8IH24bst9ik/nwpAV3h729pApsS+yTRdSm4uSR9TRtP/bOjNTtlweI4K
6j6h3Jfu9jRGGCX9IQLdlF7wqCgUPgymPNFQBImCkieqwXfVkHEN+IVE2gC6wIMH
ZEPPKOvGUIcAm/Fxd2SbAnLPlXZ68APLWTBA/PgU0e75dreeILyER4PWy7JTYJsU
oEaXFLVF3MJPCN+RJrjYPx3Armdl5+k34zOERPrl0fSwP/z0GgXJzmFJHE5eforz
3B8tZhwSvlUv41ZXNE7t6DzjVBcRbr3QmaoZ3aOtaAQFJfK+W14SYvICDqrL4bGR
hm8qblbN4gWmITZiL4dcgh3ePbby+U/mKc3TiDsBJB0WCyNZIxMfF36wl8oyYY0q
de0mjK6qjC59Lxf+RAOAI99Hjkukg9kZY0JM/QRrqRH0ChNFINsGKHBDixrE5M0x
+11VZCYneivQOvVQK34MEt9uz9AHsZNJpvA/re5nb2B+BRwX5QdK5dEvDaHfCkfM
X+CWZPCzBac2fneLHvQBlOayJW0vT7UWnjZbAkozH/9pM2NlQD/yGhMEKo277gSe
TVW4XcBSVii0GyXpZlNmqBbpZAdY678UHtbQeaWPhzvnKPF8d2OW4+TshB/ZPftG
XSafnVqZwwFQvZ5+hVXgsFdUy5xRarVkA8wy8ZEQ6+aqEGidXCBI+Fc5hX0+2XYe
agb/n3TjThTRNB7txhF3ikeYG+BjM/9Za4LA60IW6Jit6v0HOGrqfRD3Te+acgR4
HKz1Bx8AwbCNG2Krax/Yc8DZLUtuuWlxeZxPTWRtdIJuaZpQbGOtoLxO/ZBUO2j4
5RmaaHWOprIYtorcqDcuSjybcKdpCoRKpPcwN2hcdp8s28uAFQdLcqJmsjjrXn9x
IJcfFMbL4u6sH5LtXz/g60KO+2Sl4MjJ3pWJyQ1P7bUUeMD+cLKdiUcmQpmWKMPU
FKnDp5Qkc0gAAjSLAJXmxtZ1VQ1NPUiwXCjuMSnOZUIKi3/hmEPgu8wazQ1WelZY
jtm4RDMLGu9ADWJXRnXwqBdBItMYROKNwQi3KgxaIuTSOForlbGC9pcm0DK7EugF
7BqTK+9tMV4DO2LZOT7NVdCVraHBHrN6g563PzhUlMb83ZWZXUcBUt90ELeWvOzy
uV+9a/gxwc1Nh31WaUrVLTw+oiB1u/K9HAQ4CGb8KNehOuxRpM0dvbJhGDXYFVmN
6sopvjEj+H3ijkyVG4RcHxSMIpocF5eBJbUCn58iovQXIWVGFM4mH7mgE9wftoq0
UwC9P+mUxnewPUA+WX0ezhVV/7JHnw9zfKb2pRR0sXbYFo4RQumHZWE2qZAaVMRE
FAXvZGg9oleOPd6WnfitoEium5e/mhXxvxUSvMDHle3AbadBudg6EsCAxTQrR9Oy
GPGAgn4K4POiDnH0H8M2p+k5jBlCecFab26RzMUpgSby8IZRkg/8E80xts7LJtNv
i2BWvtIIq5gQRSUzEdynODKG6uZFNER5BG80I8Mb0h5jgtkjnWQzrCiL3c1jp3TJ
bacYRYZqGP+VGuPq87BhD+lNRQkuqjESg8mh2jaRJFzPwCXvvL5kZwQvaRmOpGTU
ImECkRkpL7fwR/mMkvaDh3Ta+EXRXYaJdMyMW5JgkLMQTRQ5tqYjm0R5Dfh3pUZ9
7F1DUQiGxMh9I60hxEifROHvfBfOSsm6lkQqUXZImrrVPGSjbciTfoasa9/TiIHV
wrWTzhsh+pX3oeYPrEtfWfx1wsTjjg6J4dnXgxQTkJ/99ktKcDzUgHQmmWLfwqrv
fEIuEPFDYcV+I2OggEebv6vbo7/pc64omu1BIL5KngAJ9LOWHeXH/dXxyn81zzsO
ZuKboIYdZKo3OnIqk1mRHwZV1gztehTjZ8l9tXSAnKcRJd76fMfgAzdAqaD6T0+B
5NhyfVywwrC+dBjzypV3+sKJjA+qwgPulMKCVO4gFYKd0KIbSkHs7gSElj3OGQJU
4EtZmSdjremlgaG3L/2ujRcEU/j7pc6ha82q7QPwujxnqB5nKe5Z1zg8GXRyXfnx
6YBdDcPLpuGCZEcqBnqyHFFpAFQeWbWvce/YG2miVGjNzNrV3kblqrW61tFM9Mh8
M3lIGo7WiGVQk0UjQoyWIsNOMi+XOIGfXo2DuEKtM4WC3HAI7bj32C5GKNbqapei
GBndn3pXWmBGM9h4BCEupaE5o5ANUR9/A+9ktaB6MqRTO7QTDZWb/NpORBUgze2E
UtfkTiW2d7NrMwboN0hnwI0J/+0t3cEqn/ZO4T/+7pnw7aBnDC6d6XN/IA4KJ7Wh
XwNWnpEmBa84IHk5XjztVk3I3z29+kX/nwlklqhCIagBHMBQq2tKgQbzraMw1zYF
H6VWGxR9L2+OpVpgX+SMDx+DbYPFzRLMpu38D7Lemjr5dDOuJ+l1f6bKFVbs510i
1+LHgKP+jPDkXoy/m08CQ6BLYoZY8hMRHURq2stIaRhheWXg74YlkLPt5iQOULVj
sXXdeVtUH+dc02mp59cMYgH+zLqbveR2Y/nR2t2suB7MIK+6Y+Ev2/PUUxlUAdTk
eaVW7yK6o9+SxN2ZFZW1QzgV7a8b6vuTQCuPxgkMN1xa17AmbeP7Oc5QAZqAG4Ng
rpc7/6CJsLVWW7xdoPcwpggfvD6+WtXtATVwSG9Rs+a+FD4PDm+U3o3WCJqJrOw0
dsJlddVrxr/VisijpIdT8oMbD5/oc2+EiZ3lZunftmfruXwffaxRqHqo9xCKk1i0
o18inHAgHLoKW1fxn1NPiIJ6X+cwExl5CifrWzx+n6O33RVVhxzZqOsOPjXDVR1J
0rJLIUiRTSyYEMRaprP9TPdyQc2h8rMYeMLfayl5RJFeuaua0dXwCKJWmGk2pR2v
T+bn9nB0nQCOTy/FY/W8NCoWlwyWEZaVwYt21lj+t7gpLSo8TjUBkkAB4vF6WpB2
yP7Zg6pu4xLbfaJzjsJx55g80chK3z7h6e65BalDaa5cJA3dYLtkNukU3zyiGxqm
c79ItIwEH4ysGlc1Xl8YYU11N1QtFwZP9on+z3zfjjPKS5cfdbs4T9t1HOa/SAZF
0RbAQ8HaIs8qjWkO9tlWlMYtZE1UmZGq5DCg/YVIvONn89wMkQQiYbGmsyN9UFFM
33ahucNCIKG2nKx0yfZjHj/wrVYIup8F15JIzVALTTs9QfWgaU0kW/ISILPnzYRM
mODDJqbZNestE4wJq8+V35EVZ7QevM5fEAPkgQyVWqUbfm8AQl+iUZj3mTLeR5Dk
KgvO67UKKlyFveiPxc2RyC7jnGoy/ypsqjYyYhlHdi22xEWkhxCAMwPQudfm+cJ7
f2L2KWRqp7H7geVAWMablucPO/MW1BwQQSx4lVOWOC1WnHPp1lCmayDF0wCMUFoz
fTL0WPlKx1oYQq9HNPYmvopoCclmO+Jl/HoJNn3kQsRvsLKA37wAObsKJoJV3Sj1
FKaHjraf3eRFa9frkSbqUa0CMzf9GBcm6p3KFl/KpdrAEwxM/geltx2/3acED1Q0
GvfRvZ1fAr2TGl8jCjZaP2QxXdT6nOHRvI4YPeZmug+C8DvyyBl29V8/uALMQhNr
cxeLw0hh6fUDxBNRIC06rrXWnyWija3siyV+AzlgQ4AMvgx69AHQ4meY0uUqiujx
pMpwXhgRO3cjHJA9ozGblCRO3xtlGNVgZxJuYV/n2QWtclR4UtejktxkZXsJUPhI
N25J4engyelkm68rFP9Gl3YES6uy6cTv4/1+Qvo951Gh0EtcK1oBcqGorCPIYyUE
fBVAbx/oa5yfwrrGO0tQuO8n2KhCzUNVTBdMYVumT0yhbT7SMPIGME8TIeMjWBvS
ePT8jPN04iH2Z2UK30PHaFphu2iHPNqEjBBqeXg+xlt/rRZizbCzOoTE8HOnw04q
Akd6SfGDsVn0l+RBgDi18dTc1Wozoun92yS26Zo57yqrUOoTabbKTcML2CAzpwgv
P+5O7kTh561MKquYbT3J571VPOn0gWRdX4VYL7MKpFUG8Ne1FQCi17ju21pmbxXg
VaC4Cm/5WJ7tn4ZumGs0SBEDT3L+RqM2515TPHX2c+fOjgCf4c6wcwW6wJAjTO9e
kQ8wvpKqBCa1UNuqDbQOpB7PMOuc5yNP/DuJGbzHJxXhDs7oWW66p+CuSVYMa+gs
JxHVNG6naIRMMvRFrHchOZ5mEvnV7StCBbVYx+q1VAH+Pq//na9jDARg2ks2vtVJ
he04dzQIijBYrEr6OGo/ObqKcfqlx2NSSPvT0cYv5ify2EagG1LGh0UG/heLqwAi
DUTV4qw3SAyKB6RgViJk48ytciDjDA7MnV64e3lfnmJygAx51TU/38z96PM/KAdI
0Gep+D7ZODDnZ1vdb6uoxx6llgD5keCz/p+H4bcOpVaFBb94Wwn9n9fonecSC0zh
u4nx6H91OHeVd6jGon5fjsUuQrPR54eZsJYF4N9ediiT0JrSuTedzvj+NKt/V6ZY
ANQ+9dviwX01sb81ghKp/KNZ6hucxlOIPr22+HwDwgTdIRwS8rU/X2130eAjGkB0
BaRMaGTEH4ylDPyqh2fZ3y45xfIhgcOx7yRzA1DAnvu4wmGxpgfwnbSSmEK3lgW/
KFSnvk4sRCvGMKpz+oUFujvI+PKHwiMGqt8PPULa0KVQk9zhmukG6OM570DEiG0z
ojz51JN0e8X3uwBWzNv54gGYx2sKuZZWKYsQp1ni4jJ5/sD0ByaSCUdxSHNSB6Jd
EUmQtvMh7875PEKuNtwVmPiqa4ED9bK+egsFhkf0zgHGdD4qeQJYNu8BsITRVQUA
Ezvus8DleQXkYmQqZbrtaC4wRg7LGOLyJPaqOefR1AdSIvSOgRkjDklftG77w9aL
Re8CCXTnJPxS5ax5XCW5QcApSfrd38MGxNbUvjtW5zz69sd5FT+AGP6+vSrAYTls
pgq8iB0N9IF859OIU+M2AtJhznt7pIcz+2yAiTh2e3CXjFN5KzayqVxYTL38Tv5W
JGsVEAiui7lkifLwNmjv5RVFNGlv6dXM7dBxksYFRNs3s5p9JLNy0upiUkseHrLz
hI/UuT0sMvNyfZUZ1Y7zCxMBtipoDXzKf5USLzjFiRHPT7vdipxKg9r2dmrC8HZD
4ccAutKtIgP/oLG/czsa4j2GVGQ7gbSBU66BMPP96jzNVg6CZN2fn48Fz+ZkKPJ0
jkobQ3DNT3WYSIAd0r9OhNvzIeoKHhk0rP16BmjFINQUUkVM5zvJF7DPu3GwAZ32
GPnlYW/UiS2BzJbnNLoaInUM8krbk5wLQxK4I7EaKmNJBHSjR2Rg4uE5EcP3ZLr3
VI64d1S4f7A4sQkNRVeQk416yaFa8u+m1u+6XPk3mzjlm+e8AJjSQuUSzHzgmoyD
huoScSL8ZKG4GRWPEni1WjunrTLorpspzGpY229t/cN2G9HCvu5mRdai7DLqRgvI
y+xOFysYMZTP9BF8stmgp60Vg8eYBUrEVpf3x/FoYue8BMdT+E/Yw3SWtPV9qVD3
Mzt0j4EwbbBurh8Ece9WIr2AfOw5gT1ngBffVdJPbPSX2prrtzQierix4F+Tn0zd
3FUsJdhqGlnKjSIIPHOPgfm739XbEV5DxlAv6yzzxiYmopUOeyGQ35gnBCSofkqw
ZTDfnKuMV8vVxqxAL7qHQcBnrmZoidvtPgADaCRb5/n9pkhn1j2omdUO0NS3IBF/
kobnrI9GdC6MmdkKUXo9QOsbJbDjRwb5QgfOYjHvm/+RvKkm2aRlY/XOwk/B7y3K
iiML234SmwhcpRDt+u8HAyO5rsTQZtlOmg24I9PKX5PCQAiK9uxupCbNWagBEx/r
YaPVzeG0X4yqchp4MjJY94EBDvxQDcDBtCy9OrprcFQuRyOmEqThOBqxDWjUjSRR
EJvKEsfw2/mgbDbvD6VngmzZLJAqn9EIJcmD0OIpDBclEiUMDqrIIKF+gCpZhNz7
fNseeUDlePztTe9sjujaia1e8WhQtesgXhiraFEFR3dOwb64VdocIJwcut1ePpMJ
mqSIsWlWRC9liohdAVeLHm9+kWzMwUq4YTq9z8/RXjOHDefseeYeiivoQmHlyUZh
UtTJWxEC2dfRaXFRPHgS6ilXoxCdbf6mrqSCoE2NB/r/zZrkn9Qrnfodcu64aFLE
L2ADm2UnFpQdrGdCaf1evH8SuI+zu8yG5QnkoCHolWycP/nNBfV4vxUS/EJKWgS9
H6s2y7/Xe45La5EgwwnTg8eWkAanC1uty++x+v/gxsPzgCGuKHP4y2/URu8bnyuD
QOSyUBfta2YvH1I0Y4RlB7IeKLRgh2MyBIoVp25d80is5noldWejWrij5hBkbuUK
+aviMUidyMiewshpZbq6ohMzY/ouJsn9HPbdwLHn+X6HFUL/nERPyqnY5MOJ0ZPK
JfpwGHo7y751Jl0GKl/iYUgiI/ESfv0qvP8OCtBqIQqmASQumu13BPVNLJ1reMbD
HF6VBx27Jg8mdP3Os5EiB8s20U3eJaI2cdu15IBo2pkMC0V3ZvbKD5u+DCeP2sWt
20GkOMzUmLYMn6p+Bb5hF71C4oiZSAMB5UOkmPJhwhKzSRLtgL3Wcv1Qk8VWX55H
GOz7em1q3SXp+tO5aEr7RC/9W4HAf7OvRC+KIZ6VlguXLdUfc0IVSDUMi6QdQ8iL
WjxwbvK0JJD1U/w+xdcxYJ2UJlI0WJ7NGmbyOUonN2xZRxa84wjLBgPBNOvuFhRU
7V336q3yruTIMjek8kQSjAgvKNmqO04yEhV2PihV/4vVrkFV4IgKIZ+HOwYOacWW
J+5ZyKuOpI9496yo0CUkUjupjmHB6vrr2rWyiAw8zBeWI/5/Y5rg8iu9r02t23WX
+Iys61V5IQZ8Zp1yCSpfC3ynCDuCSWemxxj5NDJAUyx6uBlc2I9qik2lAP4//jXG
l0FzRwqlV7JMpkRBr+V+IOrY68frif5yc39doibc39YXyFHK2CdNkq/yuQ65Pmap
0goeNJeDiAG2cCUB2J5I5X+dIW04S62h6UapaOw090oN4osFFiWXpnCcJ2oIxuyV
cTc9y0aMJdo34xQLSJalsqgH6cf+RYC6g+Oin8TM7PyboNTF2uyZq+kOQU/ymd8S
2xxcgnbhcpadT0jpx/6xqFJBRH8nUkUssqGpSq4wQEqjB5CavQGSiWTdJZi2ef1v
31iyWx+RVa43FErVoW1zqF8XkyrbuDSpRrEvgHJPafzDyjvumE56S1gJBJMxxrNW
5DyACbqC3cXhf3ySAZQGYz59USBrmzvcoaMDmoAEWbY5gj2tDso2x0skmjU79eyT
PwGv1Z78upjtPPuZvPX8/HdX6CwhyffCEGjPTz5diiiOJjfOxYYDB/h4mBc2nRUY
0sENRSstCpDrsUZMcu5D0oIeOXxod1sE/tCnMBEzmlN869j8TwM9YdwRj/wklcAs
/KY3oVBMLCp56Mt09wI0DSR1Eu2rD9Ec/lS+e82Gm8J/N+iLIj12+kqbUUDbtMIx
OqLIjBgoRJ6uhwoKro/B68BF+HtMz38HlterOl6l/XbIGl1z3wDVYzc2kNh5/eqT
a9DroSIHQP+wpt3HojorZ+mpfsNwKSap89DWZpnFYTmjZYQu6/meH55y/VANYVt7
+JWoBcFYyzZmwTTFHZuLGA0/6HqJqaR+DB7p4aTOcsd0Qt7kqYQivV0uspBiniN7
mov3zLDHT9Tf/niGQoDwvH0hBADMDbHO2usWApNXCMPC2tld2t9KMRrA17Ck4vid
L+gF8A6t/iKEe/S+4zrnuylf0400uFNCmMiFtJZkkpsvD6qSb0ChEvIpayGlaMVX
EWHkfSwMhd0WoL7dfrZj8F7k+WlNvNnLIowpGZ2HBfXuJtE4ZedGLvGUVJjnBBN1
0Mid0MacU6NxUc5/nBU2NBCCCpq83gaV5VjUdOz4wUG9QdOCU8O7bVWVW/YEvW9q
cq1TBTc+XejzmIQc0hPZk1Ik6W+VC5sjI0SxWBEZYPt4VZIOPuReUL+X1db6fW8W
TC0EUSNAsR7FeaDQdbyB4mHdh5T0QwlcaEuVBPaCrStOhFtKSthNrj83iYw3lIik
4vMHSU/nrtgJmxoAXEDafmeE/AP6TpVJw9OCUvchJjWZ3+UeXIY1oZ6uvq4/jXQg
DvPFTaMJFl01BrwHxESK90OrFHKtTDYnemL6zHCz4pGEvTpa88rJ3g6qFmXXZCPj
IZF2GlqcS+rH0pcotvfNH0tv3JytMa7aGOBmvAbpNe7DfM240LGAZt7OJswBSxMw
+6mfASK7iPnvHg03JiLBG7JOaDPmutEb1hikyjMNRHe7ri659tK7BF0BAANMy8p9
Py20/we4s9ezeY6Ra7y3mcZlcd7W9I8pT8/xOfbV9d/Tqeuhv3CwFxacdZSublC6
STzj1VN1VT/wFR66bEEoe9bIqVYeAsH6Mzb1Zse2HGyRyBNfy1qBzvoZT6Jsne7F
zWFTw6dP9ajDFN7LXAnmA6m4hcbarybqmqsrKuePDJZ3ph1XLtU/VJlzQZFip2iE
SFvZknk738B1sn8jKdNDVj5lQanAngGy47BMDajh8+KypnT1aD0xska5dp/mM/EM
7Hl9f+8vyOk9ApOzVlgy13hQHAj7mYh+gVB1UnkRCA0S+EF+VXeKVGq76+lFuVFD
w4NzJsBmrKETOqe3258AKJP++UEgcuiSRqJh1tGTh+WatyTKih61wVFeL5RhI1XR
HkPLN0x+zrigge6EOofkcF+voefqeFnV946HjiH7WzzwGwFWn66KkwaGfe/4JJtX
yhPDt7twLMHbRxMMnkn+ybUQygTx+wtoEoqgwg8IxzjESErhbb6zDuIrmzZo7rcN
ke36jIpGKwmQC9MelTP0m+RUv5O+0vLpeGur33jTV1dTu7D7aPxOlAKXxcan7TB0
rzY+jGBt65UazNc9S7mOZmwxS68v5ZlPSTaW/jygFt8a/APdCGT8nhJIhg2KP65N
cAWuxhZ6lKIxyoXeSeZ4/4K1wIJyoEmakSoJCuznsqiTcSUPpj4w9fnlz83nLvCZ
N6B8vbfjCi75Ii5URVQQK/qyrkuRG+9PVpQPHtrOMa/qiqxqZ7VRlXjKUyIZeNuI
f4qVoEjbI6+8ekHCVEG6OYZY5aP9Ay2YSIqXO/Xyl2YHMEdxtZocEjf14+vRmp4I
M63nic7lDHGpyojFw56pOc3ItmNVyu5WhUTmCQuWs8LbACM2rYgUyPo/D5lV9NL9
OIYB6FB/BPUkBmlPdq0JZ4fdLqFVQeAV1PZUOwFEJnXYUqr/T4jWHAH351q3RwWR
FmrKHBEvVGjjuNV3ko/oBL6B157B+tjdgJLNGCEwrvOsy4P5e/C0EyEmfgdP9VKb
wBNvE/DNGlrXDSgdog28r3Ek5VF3P9daBoa2UAvlbHattktFoysYfRYmxMigiJUd
PQX3VOwEtt9MkHGKFD3A4UFioaT5l3flA1+FePapXXS7D6PpzHyGOrA6IXnqC4Ux
wIrk3ixBt7Wmv1mb12C1wxTY+m4ZU/+eyPDebO3sGDt+zGR+YL3R86gAXVrdgqLh
nzV/xBB3tQF7MaAOkYdiKJokPVFNEcjK/HAx4eOERRs4ljwU86kqEQsOrxWQXuS/
gTb8NSnV8UGKHGe95Uo2mLkHxYc5If1U0NJ5wt3jFDtuOPvbslbLIt/hgG0y9a2j
tjJ0dyOjOgiayZxy3em7u4QCWOvLDO2gJH2tbDFvtOIE62eKHFV2XsEBIMUkeVZl
5wT6ajc0qTmREcXOw8NE/6+2kNqRJF4AvN0aufjaVp2j1hRiXmABSHL/al1/weBo
mBmVevq2RsNBFYeVarUh3rd/wcTSkcMXPldYjzIS68Pday6Kx1JPMWtwQcBEGWzk
4BGI4zXFOpYE5Ag2cqiXtrigzGNKBvhGf4o9CZoiCmZe6bKh+svqbD9zRydLCSbe
ZceIEwL3YXTMvTO5vFulvGHgTLjCz20SIJ/gkPajeNpr9KVEcqXxlfPM/Eeb0USH
kI6kzBjvOcbC3OPLPIppI8XOrNxgIFrA2NmRun0ArgD9GLPAVMrgbnPWCjek7Zlx
bWYDduM9Harp33r4WdeMib2J3M5eY7YoA4J8z+t6lG2IpgRxAXUdnvkyTzq9ic/8
RA1ezyY7n3LBF/42CQkcNU/r+vo7ftsaWO3hyu1gMVdD0S4pqAkckM1LZGV8REu2
+atOlWIE1w/IjWOfaDrDnujVY4aZ28RkbEYgDga2aPQ4gDlfuzxg5WAZThzHI8/1
/arYCK9Eq4m1hlgoEKBiQcSeuCR6i2FxtzgI76bzpkVlWbHqO+/dDMo6Q+2OXyDE
gjo2rQIJijES8QOhUhdjhaLrV2nPZIFVJl/vcmLxc3ozLkZwWKGzlpg9UkuzE1HP
cxQKIt4s2y8sohLvGPiRRTUh5WrhBjB6WUg0DQRM1nJ/AgOapgdYn78L3TIeZLsC
gY015Mb3LXyCZJQhtCxYuD4kSbVXlQg41POnZ9+A9BaRI9AlrepJ3zROQevQHyL/
jevUig6blNMbejTqfG3eis516s4wnzlI2YRK1Ojy3AEfBNFIGopB49iNAfYqHMLK
vLtOkRRylUX/Tno+lYlPubtFTNngCsgQyo74l09BhCv1XqUCTa8KgcpMV53txnsB
Um36I9zMBYgCVPle85oa/ChyiGCdvinui8a4xFmSzUfsQUHegHLRT0/j1YyCiC3m
jvamnCxP4+Z/QHaYrgwzo9y+p9obic4zZeBbzT7z0mBFWIqLXWOlM29f59HaCCWy
p9jyoJQ2nKshkMG0QjlU1nZR/zB41ld+SVOP4lFWmQtHn34EkgwrLGjbNO1AVAUw
EN6LsVOoAgZRr5FTpiRXXiIHLvajPaFXkzeePhVqlsrflII2ekntM7rK2fEoXlPx
x4/ccD+f4xWAccw46O5efUCoOqZT9r2tYtlX4EEIgXXyVRvma4bDwekWXaqhvOLF
eMpI/fmo+vEI36OUcbut+cTSrvRz9/ICguqu4FaYYjqozXiw3XaT5SuXbW1As62d
sylNA4Z9mRt/reC3tvPcI0MBw7K2Sq5qQkY6OelduYGxwgoJJN5yixXV74ktwJCx
4W2ybTRsDtAJWt++KkM4FRfw9VU3hqJjFt0OAFXcpmqT7oyRLESDoDkX3Z7EIxet
Ecfel48/wsHlB1H2Lz+fqnMOJUq0tfZWKVmgkpQUsNgJ8bz+J2ZRc8jAFx1d9Sjq
pSEF/xM6+SGrvqG+yO62UAvbaLMZ3ssC6f9VUiJbEANV62MWDHp2r86TWta1jKdF
NnNSavxR0UkdejhknFj41nqyLGQ3c7JRli1xjoAne0BKb8TpK1hGX/V1bQlUcZD2
H9EBhtNtArR2P0IqOjUs/Xn4BrkekhSapN9BeUFWUXUJIE7oH2otNhsuU8lOnyQJ
Zkt0drP67O+TnjEPxC/bIpV1T44VGTHf+l33C2/uPHxNam/UDDvkqD3wHhcCMv6u
od1+7GMu58Cm0nLX0yYM1e94mlCjtdlCnWYll3SF8iGwhM7nJ8uFygnSZV/oJ3Oz
EDUlJKw6zr9T30O2Deny1N1oP9mgx5uB9TPRzkJCQoel6dT7HyNkQcfoXFJvTskY
PY5BjDPH/lMRotYj8mPtBhQkcBBNCvj5hym8tFeYlBEvgvUVPWDMcAg4eZUp37cJ
fbSxn+6SlBJE79iargA2VdJcEDtiHzhx5QuRhLgNA/WiVg7etl/2hDmB3th15/2X
Dpfdmj0tYJr5hyZpbyk/GWEGotBA50O3e7QNiONLzBP9Q0z4dr7glcCyHrWmwAPC
sb1Iw/OyxiNhHo4fLEOJ7QFgHkIjKx9TNmSp+nXWWT7+oYyOkJUtxrjrFVKVf8S7
btv54OZs6NjHmdgOUGwZY2f6CvmCGQjCaPe17sOCttMiu1zQxT2ZSOVqzCP6fhCb
/I19x4wgLiH6HN0KaqHQNJCtHkRs5ldDrBjg1OINr/ehs95U9ZMeTLRkXwaRzawP
yzHh1i6FhYGwUFSAMcQm+j4lwFwWKbNUkr6iwfH9gOA0mXezEcblzK+qUL6kDpNH
7sDJ5NfWGAhH5h1WdOx8jblDo69mACUw55nLfaJLBxAeQFO+Eu0WBz1NpE70ZUX0
5v0yrnJEVswgWrYXDhF2a/GMiGdFtXw1R8M5OdTyaYoD9Nk6ox4rvmv9xHwT8UK9
lbt025APkMblDU10GpxjCqpDG1ioM2WPHv3XDlI94B/rp/6u+vSHRp9I6fFO6Bqb
M7GKBbWH+oBnStgSue2WZXCROtM+L+HZbto37NqAmeFBeeWi32Rg7+1bLZF76wND
dy2T0XkaszOHaLhPbusV7GGAb4wq1mLKbaOP7RzuXRTgQUlvs4wvUpjFhrsGKpNl
WvmCIoLyzA3/RfrojpX4XtDYF4W2lsOYRD8iLCvJBclU+R50rJOUeIwppLc7+dH5
vTtUSKQ+rMaHentaEheg5WstsSgHo0XTRv1uuXhLIlINJ5wlpAS+2ojt6j+X3dEe
+YCfr+m2qiVVHCfs9sZi8YQDDMIr6yjgB9CNlMqA/g6QGKZiFNxYlFq9QflJpzeX
Nb6RZbGxaow+33bqGx9MRC+0CTGUPpg2h2UITJH8jcAx4w8uvt5OZu84/6qkASyU
gMjzvqzO3nYJBoZQizCP2GD0F2f4EemageBcA7tJ2WMkDuX4i+Z4rQHJA/ZaFTtT
dnig6FS7WMCXNDykraQzEiofuxyuyrCqECX0ukrQ01K5Cey++nZAcX6byAVJIBrU
IiEn9tziETwjKZsF3yDB6OE6f5UkKY57Aulfg5sngDnZ8PB4PomJLqn0dlN1wwWu
xjXMxTFvbXUmcQLDmvvHXRYMYs5F8P6QTYByunPpQc8aswY6PGN3xgp94F4PMOwk
G0YQdu2P+7cnNGoKH7Qf7lPAygfqkorb+ZQwEcEaUfTOeAm2DsCCpELLhuRTY8HN
kFSLHAAyKziChPz/kik9SeiNXspXzOSjkVLad71pZ05nZ9QUeKogdZHiXLZgZVdL
RVYwlr+5EPMiZ/m4Q+I7TOUim88Ma+IEyrQi9UNKLtOMSDWnRaqLVwm2zjR3Qneu
Ym2PAamOMqO1UUVVv3l4MEVki5OTBEt2kq3ELSldoEisok7N/3hI0dFoU5cR8vlb
BFLUVJPJ45oTMSlDCfNlDnCSHeD+JyN64z9pNymi1EPXmTFyQ2usWPDG8Yho/5dy
gg/281kQ5ijD58HYMb/fOd/msxsVrHPh6bYOT4gGCXDVH0V3pS7AoxyLbkfi2kGK
eor4oEjx0oRObgXLZXycftpxKNNcqUwUG1CeOJtWubdG8Qo65khcxCA2ARfZp5yG
u+W3TI9YVnAdkBblan/4Vhq3be21K8Ub9jp8UsGF52z53jxp4YJ6zopAabsvrmGD
bkxnW1ex1yL8EgOrg+IaBvXeaYMJvFh5DDt1RN0b/zZ00yn2qw7DCPhQEs9IJSWQ
jdi/70VfBmpRDw4oiWyGBrLPb1kiG0kw/goqdKRIBrUhkpx2T6lG/SaPV+w29QWK
xinVCBCjdt7VTTytyCocLKsLHTwAsvt5a8iYTFVVLAQVZtCMw7RhrbFBcNcCpD/N
gQBAhmA2FL0q7G4Du+9AiLTwaPgmcJ3wZNLd4xVj7hkI5FBeNLkSnG6WiOYE3Uiy
o3k/CcBy72oRtx9xG9H5EHDVoG2jXzczrqomjhLsEwU+OmPXNVB+WSMro0vGG6Px
kaonueksC3q3+AeZ1YKruNlcD1tWMKl/Ce8ecmOASqEevE5ZFfHLZdAduQ+IloWi
xIQB53Vnb/aV2hbbDhUOAym+Lr+rDj3Hy2Qfe9ogGjC2OANkJaZ0xiX+aCZkzoCJ
X9JGwl6D3GWfdSvYZP3EgEWwCH65BJ/UytmdMIUSNdlTy6oLbBpY3uoByZiN3/Q6
PzCGmgRJ0R5or7zFrneDEzKge5kJpg5i1T1ChWx04rQr9qhsbf3k9hotoIYxKg7c
N4+OkPUULTFkz0+1MiXghbywxXpHywU3bhPw2n5RqCKgiug1oAVTrEpDT4mzz9/p
Rl2vo6xcdJn5UTI1eC/3AYexo9+L0ZGCMuS2jLJALYlJXXCVEYZtDa3PueaZTplj
5cpASRmb0npgSuqZ/Ho64qxvNoIzMaZPCmEXZK+YGEHMWKJEWyMnDg/HVYS/v5LB
K0yAbLkoMJvRHx5UwmUEFppJ4S12qk1MNwIhPFX3lfowQ5FcviosrryTXyZ+xcvD
XFZXISwpUpxycIS8nNCrpRaYvJpS+yCc0EWwCBNMaNlnBQoR6mTeqXVPQQWzkZRr
t4ePP22ej+bjd4NKjF6xUlFX3+b4Ow/nu5dj9mNgIK0MHAydP+jaGZQKpLcdQoV5
r1KJiL7FjO9Uq/jKQemxKk/qVqdqXUSFHWgagvxfTgTE5eO53FIDHkOtFm/5wPgt
bV1fLVOA/DQZpRAZ1sQE7+xIanxZGchDSHuB+0aBMGyrQOCIlW8lxBdq011ohvmC
u8gOCjUqLPv5LZ1Azu7Xay2F5jrU/xg+ycBQslFqYio5FUKgm6b8kTAXiR+5cWUB
eVvP8sKADx77gVGfVYILx2/iMLXL6SmjPQ8Gh3AimYaqlYarIAx7I7pQuHoxCv27
nVpO0PSmb7UEEs06R3FAXTVEnzC60UjqeVjYljyCiIy0a6TxmKi95KOKKQfTj11M
Q12v+T56AaxSaQuaIksq2f55pQqmIWvgw5gyLapnCJaAl4A/s4+g1gITrkwn1ma9
uDBsiBfIssq94lk1nf7iqAw3yNOvHIUdSrI1LYtyBGn/r9SSuQTCvKmxaKiBqgy0
TPgPhak4GawjFY7r4RrRsS/g0HWAZf1il1e5Td2rHbeLhFVnCpPa539zeCL7yp9h
rrQ+AuBp9b6unEtwetfKv2UsSSsFjnrzxdd9rojNkF3O0V3bsw7s9f8Uoi4xNeK4
6HP5TmYlT/jhiqFr8MQC0kO0rBHBCBuOx4FKNhUysWpoURSvRAq6yEjJ4VU6H9Dp
kjmVoe6Fi31hATxWF0+BEm9wRLtYzq2ejzQ96Qr9mJ/TD2BTnEwRO/6bglfNYpED
IFiyM6PzkD25YgusuPQp6Q383YWjYm3oGjFqivg8tI6vVKp1WiPXCgyOKxFhkYLv
sF4SkR7jkDpBSXf9MlbjhF7qOxiiSF+FJYiH2zeFVjxSqkfQ3DpVRdQt+9f2KmF0
+ng7N1vcM5+q71UJz2OB6UIAS8E49+G/xH33qH+TfmA4dKK/mLh+fFNxoCl86wHN
hqhK/Pv72AUYi4Ex2a44k0S37rkcF36r1ETybXCrqFk4t0uq1PONG/bUq2MET/uz
dWHEmkA2up0kHlAOElpSrEtoYngkF/AnguXeR0ZOennv75SeN19/cpoR9g+lGGe1
Lgl0e1g3MuQWsOk+D6RwtbEs7ZngLNQPG5mzf5RWIci0RRRzsBefGJNuLCXCMyzg
b9+KumPAkSWs5xjs+jGEYcZoK0IkHqc21cNdI/Sl2owLv7FvWEZOHuzG9En+fHiN
uIuDEbtk5aPjVzZMPsmToZM8hFKp1kTuDRCshVULMEV47S5KBsQ0nUEbKHPOuGhd
jp5vIJUpl3fm9oq2DMpAYeHQsaAfRVuwSDSLnSDiLGyWS3bP+YtjvDP9wvHNFyAG
Z1ZcS35aqnOxVQB3wE6s3OZ/2KNyh3eIg4cuBLiEZqN+z/BueVnd33xCHUUDHwGq
MED02gWOaG6J1mpDi9TvvhAXS9a27VO4NI1YAiI/AfUJN2iaMqQXoyPSGtvgPlTt
UvcvQiXNFWE/ZfoPLEC1z32f9AQHB0xmEibLAssZsQixiWWb16u0gIL8e86Y2PtW
J5ew7g5/PuuWVe5f2p7jeB2xoD1mVFM2WgJKimhOjaly3LqBoucL2CJammVWtA1x
Z5ZKtHcwCBlroNnCnmouh12zJkJIZFuoBAisIXN9LlOeeQTurvuQ8NxDhIP+TGC8
pplwk5lGBLvHfxygVhMUzAesymK+ieGviUwSEwXqH5T27M1HH9KySWMhOsHNx8dL
m71aAJaXKV5rfBlCkwc4CWL3QLuYdDvCufCHtqL79O5AVlhKrXJyA7uZzkazD6ou
sZXKvNQ5ARdW7dC+k7Tzxx+AHjKMmX+WljjXBfxe9qz07lQnZRjiEPJohgS8HtTT
mLuqgo4h68Sco03HWzoTUXor2Aa30n+1m2tibkUSxQ49DKizFpgbjKCBE1ZL/HEp
uBUgmdBao2YFPaq+QyDvMot/wN+JjGdGoz7Zv+b0122jlfZxo43cams4bSH+QgQc
EX5+4bPYSw8xbHqFU6zgN7ZBgppHDCauLbJ/QMl+xjY5oKQQq7MqeJ3YGPpbWEam
TD2yj7pe/qTixTvZ0IHw+o3HR4p6U76CfpBtvBiARuEjyK4C2M//fAWa0ufM99DX
ZmjUwO3Wo2R/aKSh2hxcKa34j9ICThrSUT3lZOITsjfgo5Mi0tHlaRQJnp8GCiut
j1tE5iPyKUyfOpoX0oogAomBDETIOf3HGqAUIoUlnGyOUEmERetgkTuYSEmMRza8
HqXMuchl5yilzkAHczV4NSycoSTvLnpIz8To6nr7WAHqmKSekJJR3g/YJdRDzJ32
bzguD5+A15XwzzOLpjWodFncc9Qq/P3w1VXlY0bNg4nVEs6qhadDXQNAEtWBWmHm
mQADD9gkGdDlXS2LHh59BBT95rQ1TLyVPQ7lDsirGFb1kbn7y6YdOrdMXI8lwUcc
NG1uFlXJgRr/IsEqEjEfev1jTU8PaK02yRHjlCCtfmxZYkl6W0/PtkGGw/JIGTL4
P3B7FvtsC+5rlVEROIDGfjz0oYKYvCruOcKSl6xlJKj0FHGT3jIC/EY9IuaJBoHY
NiWvDfnZ3GKONfxxNlH0ughOzISEcSJdQT9BZ2xROhhrxTHZ4E3L8UX+aVOPYwVZ
NuuHzzdwRablkzkZ9bGxaqH7cCerlDZw4ulPITqzY+PcoJJgoPo8l4p45Oped2/7
Ws0Fkzt6LawL1zrGhh0CnU6k829lZ5QGJnSAsNiVfKYhdQEmR3p+PMzQDtgHUj8Z
j8/gKqlYOwsGaLKfkK0uxRm3TPdsAFwUwdITOvuCYQUpC70TBXTbyu099l2uF5tJ
j/1/0rf2+0GiyV4TCjaYWGhuEWbrAhWJYHM10tCBZOWOrXXceyLJgBzyiM9HdKUH
R+IY1Klp16t3WWdBJgjnJw/O7WFdGtjc23FYyYDP1AJU1vJYQs8BRjRI1QD0nMAY
uIHrpJe251K0BSxMaCQjWm01JW9WNKxp2sLPPHYLrD01VFLNn+tlO4drnNdjaYUy
SwK3FSmpB8Zx57C9vgERqW42oS8GvE7ZgYLLDS1MuflSmHU4PuN0AK8BQi11zbmA
GlbQsJhn1x6r39Tkf5n36rpNG8OUhMQUZ7F2TrUMLDQUMdLQdLhuHINTb1M986mS
peoebO39ZjijXA2dDkbbFMzk2kXlcewV+xC2ZB3GC7OUSSjgecGkS5tPa56OwV4y
PKYPmhOht5oRQBJaLsA+1pdr8ufeqTwznlJ2lalhCnoy9h2BrW7NXOG66sN/aNSS
kg/u8MZPSQ2ZZ9HnuGoNY9/Kfew3iugdOLznrdleNUru1Cq8lm3h8r2CzjDIXQVW
yME6wV2QgfD6BWZ6nPYzFm9s86CRSJHAdcqycOomo3YBhiWJEYfQoKp7GOo+2L59
O9FojMMj2H5gKRxWk3u/L16qW97OIo6U1fA3HixiVFBpd4AoyvawFdW13Z9xswjf
rW++MRx7DilCyV/jVo5Pa19goEQUy3JakpV2r98JANGcHvP6xI/z7Cg3ObcGQilF
fNY+oqXF8bdaUsivHvo4pp6jhD4d8+ydlnlfb56djWGSM694H8PT68akbaRmbb1h
aX/+LZkueYv1un6WIxjjlKzwavvxPH1s90XRYROJY6/KWMMj7wC3Jr5C0JTDu1dV
e5RXE4MUZ229qP46GqMdpLN3FviHsEze08+uc4+6sAgph7ZdkfnMlG49VSkaT8LO
IFsZ05aU7B3byBrp/F/omzliv24Pxvs/j8pfKaiBQ90MnANKMPN1Y3NDEwH3UHuv
uRQw4HOihR2Niw469hrhYYPEj7ZBgfiF7QyFG3pFNHdGh6/Ur1NpQb2Ed0UQ0zSu
z5OOPXJfqIhnU7O829rt5QrgZPZhrbCijZOA9D9CUOy2tf17cl6LGGRNXVFSg+El
k6icMI+1RdAScApVKNyIPKM37m+xvTkYR+xzSUssfEPDlAC0fbj8LeKoyUhlM/3i
ig32DJX8jkIv/4eJs0ilUorpr0F3zjLlql7fXjqEZrcLoy9mfi5zNRJy7V5PSMBJ
wB90VJ0aigHzQUAf6fNS7uV+9ZvP6ovxj5cHNWr6fh9DGnLKZbu/M+Nc69DSBR5V
H9qZ9BN9/CMFmumETxMQ2iYntOJ+yVNcXi1LUQKxfdqZm5DsmuI4xu8HK4PwsJER
bwl8aimwUwt0MvGghpp1uvkjun6zvqOLFLf1EmiyB2VUHvLWeZdNyR8ywYHGusEI
4YXixc60Eq17MHkJFVGJNOrxHzAYPTuIxXfK04mWjwo5rt49ujsutPgUaliOIGZd
Ir/TM68CNt1i6s6611ONgc+UUFjChEsMOt/Jubt543p1LD357IECxTZ8TCkQAOmJ
WJ7KAS8dgo9GGgielazdPvgZMnuzeVhYC04fQJzjORrGD2PbSLFwwPQxvpVFlpmV
Pd8obxQOyGL/CpmiAVQFn3Krm1a4hOXV1lnydQKc+iTo4Wr13RgODIL7BjeCTDK4
6bEPPDuxI8y0l/WVQqKKCK+fY2HeuOucsi6Xa9/FZ6/oQt8Gxd8fiYqpMCv/5fCt
C8eNLtps1rtfaIpOSsZs85+Uasggd4x6WshPALfzH3mXeK9u2HqfmTYdmZDi9VYT
z7+1vrwViyEgCC7SaxgB2vgJ8B5BGjWneufYRCOtTkS6/tVPWDewiteq6fietQcV
ezLyuMSC7CyibUHO3XM/f7sSRb0fIzooltjcfwkFWErlxSvGL7RcTisOWtCegd28
dTBRCJjwMDzFp3QxT7DK2e0k7vCXjusfEXbUi9gjw85MQDWfpgF1R9K+u4hPL0jC
OLAyVE5ZxDPAxZQI793KPabbBTg0jDIj+QKwNFpn0dI37E6ydLkRuJ2Y59dTtfLc
ZZcdDCwNLFKuGbnw4/t4U1ykN9WaybP7iz6WhM5HPhr/kt+wTEFY8OQDQIg/oJZD
VAP8vZ6uh3P+3cg1OAWTuf/3mB+4xwPDZtGmXHzGaadUjggRPSwA9EpBpNAlI8pT
pB13n3Kf3CCI31D4BndxRHXC1oj/e5czV22U67WzNWzA84mHHvINnHbZBoPTxjvV
0tEU6Md/ho3soCxlGfIIlY1MQs2elZxMaHcwfTjQEBVXWcSah34dX3VwOWR9o17E
TBwhrVSTUYYoYxLKz3TyG9lKv5KaJTIUuQ6HXgbGb99p3Ha+j/JlJEE3XXKRLh7i
5fzIWrr4O5kUT5+CpW4v2UoAJvOgAohQeHMVhmyVVLnD21xGsFVoLanEjU2QfLzv
qhMj1bLlwVTZzSmCKUPnltLxzmYHyLT0FkQMDXm/enaX7DNQy7lfCVbnYApFq8PO
fV/Z2pAP6DmBsbOHe51p+XHZlf/l26Lbamk54DxGq9IsEiVVB+zFVyI3BvMW6VbO
cfA3t13Mb+ysYb8lPNtVN6WSaIcYc98Lc147e1mlF1J6m2RXV+LzEIVoKhBu2ney
F1VX6xVAtvJzq5XXeMCFgBTBYFeyQOoyCU8r0VC8gPCJCTaSIni2HbslncoIk2yz
GG+fuaX/sYMTdjEzi2W/gomsRLdqmoII8Mw1EtQ4Zq33mxWmNYVYUct8KLDYbbXZ
GxMCJCac/m77jAOgYd9oUTCeukqRq+T8gLsdJy7msYs+w04Jy2m5gp2CK14VGoay
J2fPz3EBnFG73izeJzLDsqOnnhDHy6wN0p9hcLnRRYq/vIIofrh/oqfHY0iIAKIh
3dIlDcBWHXeQ8bP0xQZyeb0M4Ti4yciKnUz5i3t3mqZNzBhI4ftOsQ/IXDaE8cYb
kqy0SlO9Fc1VgcnHuhndXlgfOWpqhASQ/jJI3fC4U36Rg5olUUf1Nt9U4hsIFrRN
7s1uSpdLh42kXj1sE0tUgpyeoJI6gaZubO8WEUvoDDU0I7JC28/S1B7s/PO90qa3
Dfxcm+t3KVLi38IstnRLApoDrU95bPgNOSpxoPR59sRBfGNPbAYTl5G8q2bX/mft
VOXcdvY7yrzVz8ZlL1mDur9Jh8cAikbpvJf7D0NXgEfEZuq+OKSzAvWNy0scpJho
pMUeQg51pokBxNEWGcRFHB35uDmUBcQmWiHq+eSHoojup6+5HTkyIfKkVM0AJ/c8
j4ej/Po7DdYFrQvMGbfE2Zrk/TaEaAyQQfybxAw2VaVALuyKKSyC6+Qk4Ok8FBAI
f64a/+1S/h0Ay2BkG2ENpCfdVHcFatkHub7neu/lRAJ1WzDQlfrIdZJFc+D5JmSR
kPOmItMYgFkATJZVnLbYfEYKHnaKXTK4FqSMqh/Uac0gfOj6QIv2Gu4WHVr+g0NW
MjkWszcVvSB8z4LF88Whq1cl6Jse3KE/aPUvKd3qRqNWPxokdCEtMfB3xslnyJaW
1qlnuhzhUTYytUkQktLYZTVmKAMcC3rl6JY0QGQoWTUdenvUgtKBtiL58VfbQvvD
odSrGrCExfUVoWXy+Hy33xWY7DsmUJ5TwPl7y9hjby5TvyDU23GnzyHz6u1J28/T
r9GImgO0zQaPElsl4oH48+olhI8xiMTdVzSWG71Sk4wkBg9x5EJ4HTAHI/srkUdV
I7lBMOubVEnt4xoUZ1RuHhbOvx3LSQ0X5yxOaNj0rRjtqNlamGTmKbZ4pHE5xnjs
YRvq69mvMSifz0pY4v6soyqGIyMlilgmTK2j0cDITJ8ZpbklwmmQTYup4Tgn6Agn
Iygiy4AuLdf8S6WsjucsGtdwf8a4/hKAHucQTMJlv4pISgRCt5y/nz0zwGvWx1uN
q7gQE8TxhlZTbMRlUNHW7L0N1jLFj/Au0HIWLixUcHmopcmsnWCzuQrs9uTFa71n
h9tMhSvEHORvk/g8TMwOQN4dkG72fgd87hWcRfUTav4yVgs92/QVaiEoeeuZuYzP
cI1cUp7YEfHMlwwemMgMvOK3IeHmheqZQIdeO8bUwB0ADMpnVTctds5R9NlPvIif
SHtVuKftUcFhL+vn2I7b79+AkaAKBos7CdIS9cI5tFMBs3b5xyNAcMoQO5AxbkKT
zokoWF2u6NJ09KzGytXSgn/rCHK7GvImhIu0XUdfEChstWd2feturulyGzoSZK8F
6E4Q7NnBellbTmG3YncqKZ/fSpGH121szk21DhlY6EMDHbDFskiaJ3owCEBlzQD1
Gl0iz5TwM4V24qDDSx5n3WBQOu6dXN1CsY2G+uZ/VTrMBz1HJp6NbDWNmZr8/ifi
gz1IToXWMXK3Mj1wcv6buYbYpSee9q9n5Zr3Gt4XkcZJkMpfEhGIigrgODBEZXF6
4eRPvZgA9IpDJV2mu9O2fPvF6Zd4woeVg+WHi1dKuMJbqYlORyoVxt3rbsjEbKLs
V62tlgTvg17tPsH5BqP5Xc/JM0DKwqfJaTdwSpGsOcWzKG2X0N8YpsdaGX1ukK2v
MfMKtfXT2cGrQ38yDXKgvUG0Jo2Fk6aCr/PHHxDay2hRd4L26flYrn0Lmyv3D1yr
fweU0ZjOr6caoqaJRcaUbhMQMqGALq2q3+/wEIVdXIDWBsepBoUn1NqIWT5PnZqq
73261PUCq8OqoOPx0qFo/XFsjXp5JnFZ2SOe4VgeoTZKu0yi/WPXMU5rhigMHdxH
dpcjSgHHC5RONj7oLISsU7g1pYBRg+xaw9nPeIidtwPIRnmy4dfYxKnV2gGHcQwe
aGOMpyZGadPFslokzPKcMXzUToNjwkD6DZE+Z+d8PfxVLOWySl+d4aut/uzHwAiX
ghvc7HYfMzKP9gryU5iXixR01tiAjCMJplXNaV7QfOlGViAWFNieW5n3yjPr40xF
++9QoILVnjnZlKZ+8XkFWD5lUngSApjgJX1ugu1b7pDpEBjOW+N2z/vryM6lMEr7
VrLr11Ot23PU2eIwKJQl2GI/WNoi3X3J0Ghg+Cu4yOSCCmMO6AjPscJTiUHAfsXT
LO3EZhbtMW11b9nD/YuEbox0FBC7VkLUG9scXXlATIgFaoIv8CY5w3zwlp2VvyJQ
U9EwxDAXs02CZER6no05oO7UFMlEySiYF8HoAklss5Bf6MPLYDnKY6G5s8WDcS26
9OwBw5WgHVZiP/g37sMBeq5vpRJrVHh7jkVunRPh6657grv6JkJBslV0hDxIleoL
C6iv7urYjYWgCnxyLcV3ihU3Ia/btaOwM6SpFXxKtVduIexcSCpJSvTLI9NAxz1R
dhEm7cXdm+4IR9qjJO7ebmzHm8ej1bIAJm+8dADdFjz68oLr7BwyBsVGCHa/KpM2
tWFXL7V5vcXfHyPAYl1aZqpPFvhhCz3UARlJnPhL1HWbVh7AGF+RJ8n7yvYWuLVI
RCtXCmS6uZuAXy9Z6jnGTx1px2WaEBc9nj0ywtVSPGzu4GaJolpxH4hFwBAIQZsi
rIDQFld/sNERrqoLtfwoYU/cyGnQZkBH15XSqP+oASWOjD7PlLGppsdryZ6yWb5B
qjy0HO8hp8fIJQobt4enSFmVHiouee9S4UBji09FquCUkbHlFrzgJUlowW5gOMxA
GIIsI3oWUaG9hPOr9uHZUmI9AjdQTlULr/FRetIeKB90bE7FwznTMC8Pzg7yvukc
wX/rVE0ySFdnSFXjV+vfBZlf4G7HMjsZyouIlUF1a5o0sk660iWm893j93HxdjIT
OsOYY2mLYxDZ4cQU6wrd4E8zQLulx644mtZiqfRtYdWTLsaqJT7JLSQBphjM4fvb
rcRCWeBIMqt0WUSeDsS9E1JHWUJE+nqXi8ORpZPEo2S3V/Nyw0yTEJuH0AsdU9qk
0+11Dfk3b8ugr37fM7/1gcvBeiiUicnf9vWqGqU9KHwHBtYxop15GNLzvKfdkJBW
zx6bnZmeRPJ8QXRH/UYMIyBIOguy0ZXRRGdPM9bhbyp/mDbkPvb8xiomDrTNsZ7e
a2HdVLN/GRV9oMvqiT5dzcFI4WZVU9bJy2bZ/jNMLndzuKUuMK0RHyVJBy9I5VCT
j1ZkJHoDwBPZilJuNcmXti9BUHBCSAPsKvHvonfibr8Ki63umTv6Tso8yYdQ5sxH
EsCICPBDrMJRyPqiWQgxWkcw0yhhMSpRgc8yleO3G1l5N7pDi6cgGcCUqlNNDmkm
YGnWi3uVSnVbUspjUSBXszMqiECKhVbTAKPPT5xqb5b990D/4WZXtjqdlST1C+WO
6L7Pls1jhUgMxZFwisr8Kda4wu2EXauGJTzysESZ/avtNHoAlbQ1iDNGBWt4JQl2
hOTyUR+XjNEhr7rIvtJnamqU6dHg4cZJy6ZiYUuU/c0H3/ywIxxvvb5sXesX5lcT
r97TaN6xDQPD6dK/qazcdmQUKKU8vrdERwYdWTCcWpe47/bzZKCBMNGHGzThRCm0
zL6cdsT+gFqPJs39FMp4VGkHLfFPzhcUTwWMFxOSsnr7Dk7XLV24A91NWhdAF5NU
CIk/KeDDptWNXA/TEcgE16+KcduYGxK1jQwgZ80UiUk8p5MHPI++1QgB5hQK51hj
jIiyM1ICr03FiQIpEaZxEqIPZPRMyf1psLF7MI2jYgLNLUkJj1tSS3svR1+f8J1e
n02pkLi5lIoPYFT6FEyIHxh9JeS7aOw/Pf5sZX/JT00znwY2he6RBx0Ff3hXyonp
j8K3yWizNxmuDtCJ5lX0WuWA0AWZRk/4W3D6L8FYFZLE39LH/k1ci2036srdCftT
RuA4+8Cc/rRUHENzBX0XnPwpcZXYd+YhL8sglz3SIfTjPnnXhTk0Il8TKlN4eZbk
4pNfy4OrF0DRvyNWL7demiUspCJR2u+hfpwAwrKNXO4BJ8ixwvZLTvQ+uhIk2Iry
NtT2aczyGagDp16CfqEKnAvsqjVs3Cksl4iNXLAjv58fAVS9AJCgvktPVxaw4JGm
cgaiOuDmwizaP62ZCVhvOFVI+xChpKOZAiAF0SuHPAa0Z9+uhI+rap6lUNuW+iWb
hMq/ASiINHhr0pHQSTZlCBO72eyMRz/VIZVfrnYkEIcnUIxr0KIqoMt2dY4r0rFv
wrLC8XNc76gUoEHzWsr6xT60QAgofCcT/a71kTbaF31Qx+7uDgZd+g9Nng3Kq7sT
DpAXsoMUCUZU/dVSSDo/0CmOcqjBnO5F1shXLqNjigb0Wkbw3X1TNeELcz81HFxc
Cbq2iEmGAK1F0ta6JEmTNfqvv7BCXqIBhMMRIHdUOLZTdiMo8Y5yfs1zebOeiFat
zsmWd2sU5TyMSCzwiV1/SKbGs7yzME64JJpmfqrXmdmJqGujRw5LDjht3HIEPrxB
Tpk53EQL68krGh29pCj8n4GdgaNmhfOkR1TgsqyntE4cX5dP0CG9sDNulx5ikuJk
IWs2BZF5MARnQIX01GdiDqNXevduEGKyyJIqCB0Bj4fSzopJRebDt0upq+sTQTwd
SA8oldrT7pjGOZJab5oRTfQDMbUHz89YDPEYUyKxI0qD6THKui61Wyl0AhyB00mA
ljyDETR9wfBqw+bKfAd7CKwpnZTr/eVWTYYGm4hz0+kmhgE6flU82oSpvMDMSoeA
fiKaQs+TD+37KhQvU1H2KtwMlnUYR7eTiv387+2hH7j+AtnSdUJ2A2pf+E5/RtAL
JuBU7clwU73yM5eBnAkuNDawq6uVvkoKVDyVeGYfV9GnRKuyV/nAHZK/HgKnZzhm
cwEyaM4iIJhaqddRJYuQDSoe1vTkFuA8bN0kuUXf+SZ7GxwcZSYmm+dAtweUpqeY
EGOng+gaYtJpQF6FunKiL0H/rTE9hDdjN9A6kI+4mRSrQCd2XcHrQZrIwnntqrt/
JIGAcyYQaGjsTIXp9kFtX/8ut3ThjvF85SaPWOdYZJBO5p+Mzqy0CVFSbqO+NW5/
cyWhCMFcEipWGcy/WtaTNKfxll9xsjuG7V14p56LdbIJyK9OQtEHfv3yA7yz4brh
uxs47/Wz+EGw5NZwujQSjA5cQWzcNvG42uEbAA43ibpUQsq3BsXskAIA0TUZReWJ
9XCYAdv7QLPuQdGPuZ6h3nFv/LKbs7BYrmRn38VNKwDPaxQ0+WMzwOl3hbJYnHAV
BdPhfYzHsMCCE+mCCk1+Ku+559J1pctWHznwsAE5Ulc59pWr2k9LBKfIPuyOSK3O
Jl3qvnC1TSp6HnHOTuNVbyjRYBkgMFLp94qJo8bSWyFh9eLvlItbBXR/dkGraWXC
emahjpZatP5MhZLaTSRW8nOkfyZTCepOHPPgFolEA3WChmdwkigq9Ua/T9sX9r3v
u8sesnXiU0jYcsMBKu2zdtqDx+iyLqmKF0P0bY1+HVN5TiDhw0hhLsF7FbcAGXOR
+L2lw0ftTl1Mklaoc9mEQZfuO8sbIEgiKvHl/K6tnWEgu8gYwveettw0sKcoqyWv
4HC6jjehOd8YH2derjpqKd+PzJsDkpzK56pNhoPyiDbIkybRgccSXbu+TQ9DAHqs
XwoOEyYobwmqww0nf310zAC1PoQQrAXqN+vdWzg6jTaYaF8YzTIY/9eCKKPibvZn
F7TeM77SAa+SM5jMBAALsRxkGmo9eIXJxTC6BX9zewI+mC+JXlI4F3frpWb3OUxq
GnH4Dpx0uCgXKACuUecjbw1HU3lM3m5Ou/hUhjAnw2+SaYq6auftOGtg5fAYAbgo
OPH4eRQmpNyhJMJK+PLTac72i3SnTsJ2h/H7KZWPrbrfY8UIRyw4/AqYbRYYq151
V72mn38iRVAHB+i9GMJ1UIMaW+d/hIWWX6DJHw5NNd4tiWxeMQ7RYMquMQEawKDA
Mzw9xxX/WKP6XfesEEd0qOhx4d3XJKn5AvvkgpeHchjWrOEH3un39IwrksIz1bi6
iR4E0WeX5nRwsIrNNd7xmqHtU3N/hrahLRx88O072CCsILk5WrkS/xTQQsOzcCqU
U0+yu7eu13TVRqSH58Y1XX7/Jt2GuImZV4uAFxrK+EaA4A6lQKzVgZnAeItD7itS
4v3y2t6d5lMaKcVdMhVXuisPujtOvAIEl5qXN5C+GpGPyONMhP6aYU8n3iCrEEPl
qhVZ9f4F4jldObHGCY1NI2HhX77+6u0770p+8ktHzwjHmlcX/OkrBA5TdYTkn1bR
p4767/PxNBqZ8eZiWHic+zvnNwYEFIiO3fSHUMJHAX0NYzaeaLwHfxXedePoi0fU
dFNTYjvhazY5U4DJi0uZCOMpTxdWhQ4uzlvlyZr+CRwWpNjUxt8h5FDovmgwlsrF
JH2BxKPMOEvdwrwesw2ww5ATq9r940dtDGtXzX8BLt3RThlmaY7YwmPsXxCUO5ri
EOTqHo/hmB7VEFXJxalkUnjXMVfEMrx5QQEb6F5pmPpcFnTVoGS6BGKLwBSXx7Px
GInSZ4uu9trGQheUdoAlfQjhNuv2IfVFegBM6tT76m3UZERZe+hPWnobGTtYzKRd
1MFi0HtzYXDF5UW40dll0I9hfjSXJIsPSgTxrPU1u458LoeB+R+G0os4GmYi74bE
lLhxa2WqcxV5DZBZUDO1D1xPyKpwupj2E18GGs++v7YbjLqtCBmaMpEJQCnZ0Eab
aGi38XR5GGyeI6ZEcmY00JwhW5LavyD+X9p8IVF3Uj7YoAffCwyotw2ZVUvdJz6N
0v609XKi5wuIH7pqHU3lOucG43NzmVCKO7pxlSQvOrsuaFSh3x6jJVihU6a3IiYj
6v2f1HteMEyLsao/1+JvKlmmWKuTtitQgBJ1fIFqvvzqi9xqzuBsNF2Hkvcq03g0
7gT1WQMjTgO7/K5o3AQwxpIiC37FTl0M9q6+CD5PEhELNkOOSECDoS7LU/hhStG1
ALHueQCwHcs0mtvL6krWshvYhYma1hPIbx8vqfug9OGCy0sGa5QG88SSLVZrazKZ
uqIiYTpPSQelbG6Wtf3aoMfYOvyeCcGG3mKuCo1p7xpwTs+U3vQpo9DbMmzaTWmB
KEAP3GpMn6J8Fyxq1KA8TVAkqpNvDKxYvs+a2IH5IpxfwY0gjNIHlWIedYuEnYnq
H4C+2wPDbCF57kcEXLS8E7r1Knb7ejQUx57T2vIzYxGXcUl1rPcLg/7uuune63og
9rfPpV0DaChQFJw89NHJSgBaYPAk4E+QEnYvqgyB+qXYy65kUApq5DZVWFu4mNYw
AqrEr8qjTo6EygEpA4DFibngbuMUiIX1r0N9JjNVJMwK/kXHI68DvR7zf8+G6s/k
DlmeSmklvXqV59U8fyNkoOWDH2p+IucKjnzKZ2jH+pUK/cEiZYW/hB7W3u0skazG
KfZqGF9jzPKP1oP9zylUxqqhfbsDNyfbOmsO200ZPYk7/XVwKrhgDhBsl+kLumcl
aMwZikigsnj/GSBIh2l3Rsz02rTiXD8e3iqERPoye38rmQOko6/T7MAoadmmv/ci
+4pL5Sl9LOZ/2UAtiDrn6/gvp/34Tfou8YxQXApz1GshIiTxdldu3vGpxeLKPcNU
X1IghdFnwry1SVIjav8/EKS7U3wlEVJXJlTJJwABAK9VqsXrb45jXaITHbJpfPyY
3AZDr7h9NBemESD4AQHCG3ebPu/zyTYQTUY6KN8X9hDRAqbhsVyyD3/Gd+C8TkMO
5S/Pq3QHBLMpMRXkJtpzlBCUgg5IvbvvX8/L7zW38N79zcBidVbjXudpRWTMSKYv
FaqwY7TTqmT+L6fCg6H76xPktzm+PpDwPzAnMK/YUBZilO1B9rzMZnK2HCk44i6S
ejW+IfQjXiWkg9WA425PUMox7HSDwwbqEycVnVdOnB7vM6+JjJXPqcZx50LtpBk5
Oh4AFSw+TMnkqu0fS/aYcDXNNlSygajvXBMGvRlGmRQ29BTnysd56VVSuHnOBX9R
Lw1/fWCIvhtp1zWYDSIUTwIpz/crR12DEnyUBlOzzp0vqlYUl6/RuSxzqnvW7pjI
FFTKKmnZGJTs4Oq066XVUPPqOTvMw+2roks64JaZn2ZKAPris6QJbtrbynrODRXL
m26AlooeUB+VJ5onfR1NmlAcfZWbpJVyvJ+NjFx9edxDz+2jFDB49kO/MNeRV9Sx
AQXmHlcHcOrOvnIHVuhwYuyViWzM3E7RX+v+rlaSW8pR+CFFEg07kMNey8+Fl9FF
kKYhnt/CIgjzBchr23zuTEgZFk3KzrsLno4XNWwvqA0oGCqzZpqWWOeyOtwht461
optwooguNRUKdf+zmdd5R+IqkXsULP49Kdvu1ICA5PHFIkyRV4eW0IPgft34ZdU5
4csVzdekUyVTc/w1db4dtCw+wKgwJebQ+Tf7F8XJvZGl83EXeFbine6hobeaA08g
sFBR//Q9bq/zfG6aHSsgdtjKP1NvhDsMlKIeyVSp8dj6wEmd0a1YuzRePkspEJ/u
nfffsPrt20pUD2aNwevuD+QwWFYts9OUpqYkazcIb+fiBcycJMYLf+iFsLANkH+4
kHE4SAdJVQWfvg83sP6wGinTrGbfm9t0QB6qE2s0k52tXYITgprGE0kmYJNp/Pi4
iRXa2d/cTlRTDMgLlDV36mQeeN41JQtKH/QG9Kie1GunHnKg+CJXD/jNuR2JgSvI
qvaW2n2nsJ1VsefagUkMlBeiJjd0F48PlIZfL/YMv+f3mR0GlvYsE9ZHRjIWFUxm
DB/UkoSR9Jp8oYH1GRxUEmKD4BZY+7wmzoEUXCrIqhl9DEDbgDmX41jSlv85Ffqj
0vLAPfToOF5M6O67k39YWwRRc0/1MV1oeJbIUwL/X4v/dNM9GP1O6LGj35n//2Rl
/sBxamglByJxOCmnsKD313VHS2IqbwQW4J1zYVyfYjmEdltSgAFZG6VeW2DAXunQ
bTE1d9qH730E4U4zOg9FXpbI1mrZ3G8pMADDRKc8AU8UIlXaLl0qPY50sq6T3yug
U/L12ytxGSrddPFFtPSt4yVFyp0RKzsRHnKVcupH2KAI4l80t31bZ5Ea6uLrGBtp
+X+6L6vzQu8qL2FGgsHMt+kfqXPXX9fdLjurqfKTbJru6Z2tOh/PoZif1SlMN/wk
iU4vfHutrOaCyZKiAeo0INUjUxpdGQe2wwU3xR8dpb+ee8v3niWLQK480vq7h7B3
fn3CMhKXhUxGrFLp9sIIeKe4K2jxowkW0UYIVigCkaoMK1te6VfubXVrRN1shkcg
+W/RzhhP/pE+J6bzXkOohBak6sG/2GVOO6x7EGK589BR6jvteLcWrXigAbZAWCkn
9WxRr58ZH4lJsDVRT4as7gygPt2K7qDUCn33ALSqTy6/y7IsBPIOub0tjevWNxD4
pozOCRbSHS3FPyupCpTplSfA/icOZANVJ8KkD4CUcD2PNj48i6+bpMMO2d3sGCJr
YEzKWl9+NO2VDQCgUxcW7VQ0LxhAK7ghRCHD2kOjHXzUx65KPQn6Y24zTg66mbLv
4GJ9B3UcRmZXiYxs0Rj1IcwPbxblPuWD6/VYmWp6jrPfQ0tCK4z5oEfRlbZS76LO
brd1BotpDhInWfFFDi1N8gwqJV+z1YKfcmogaKfFnQ/mYD+cnOa/VKm6oMU8DRLh
AOHpmKYcd7taxFqRewllW06G44gq1Z2Fw/ATDtMC21QpjMOxnuqDhTdQcV/XYCMX
htdIaLwr8oVisf+e0NJ60FfMVIs3r5y7NSW7KLh6HOFqqqGJLYaSS+mE+8uFJwqi
BSsdOwieCRkMif9ghGQRpvZmT6fuKN2rUamhiiahYJ+x3HNTRIsJ4hxMVmcfo/PT
AYBpJIh51gUlByTppEzY81ono1PpXEypHS3zBZvu/KhKN8uDtBFVV+6qukgISWNF
/GtuWRYwsvPCECiyh7fW8ARITM5IkZsH4jznJ+rtVz7vI0bxt7pWESC/SbSlaj3Y
a46+3KCJ8XxcYawOP/VXlnPUcWh3O7qUd6/aQ/BTOt9AiokCRLQelQnUSgfYFSiB
R5CEbXFkaSNhpYN0PCIlhD+h0EzJQGoPkA+/qzEWF7Sqfhxpotfa3iPmpfiIo2zX
6SMcARZ0258iVA/G52SBY0r/PMOtP/NrY6HQQrOkwmJc+UenaBDUclHpei6tEqUC
yRwSCe6hXDTq9X4zY3r8G+s/yAN881Wp+W3Y4GlV5nRFK8aN2UP7HV+hkKpjYgCC
OP9czGjiSb9fbbvsLjpQBhLPUVnuW+zoqghvFbM82+xPImhszNVc287xucCmj2lO
rSCLVjHacORZRrHvrnd4DzPfdKUr+4seAjDy5RWlLg6EGZ3+GdDBVyfPuJARkIwM
cPZ/y5iZLfQqKU5WHepuD+IxM0egnCCHQfJisCElqIH0gYR2zRInQECvud/GL0y9
VRa8zpX428ogqnXtw0uZUEXnA2q4L9oYM8xxux7jhJHw7J6LOYhipaXy+dX9ldVS
5gDRCloUxrtnBuRWwhKtSxLWhhpHmq3AACwQulk4/oavz3myRxyLU3NLXv1ras/i
EKHJ9AWOejVdvZFjaJQ3d3HGlwh6qp62grro7chrJZXM6EDrTP4dxP4CzCliokRc
PROTVQfs90BZI7MYl3Aqv1HBn4bR6062SGUQqjHdIi1AzcMH4G4vehsGOMjMx3JM
9JkmeX2IxrnbSS7VB7loEl0F8fsVMIASfg51Qb/IqHGv9ZJSiJ3euJA4tGMiRSfs
DRUI4KtvVIWwmIyUCF/imV2oPvYTmajcNrQXMkpJwwBnwKN/hS3UwtyMEcQf8Kog
Q1Z0/h3W2dNR3fHZVN6BU+3irZunhfcrUNFUaTLx3mBnoKXxXSXDN4TZMe2eA+rc
ITP7YcrQJDBMVSnNaNZWO5X1hGtbDXNMNbIRJ6cVEUfQAtt9MMyCozSTmpKE2pSH
eVtd2VgHZsOw2KV1iYB8FXMLvgK1bKEsgEuWqF9IER/LPyP/IOtK+n25C1I9Wu2y
QnYMTRHmyf4q/mr1n64rOVH4LE5Yv+pLfw1X3OPkTpYjw9K2xku6RQe+UeJzUaUQ
cFdvQw7vxWzhSWwVKrenvBSnC32cG6PjbbGyjtJk0JWQ0aaeahdzh8X0mO2QA/bV
Spunoxebz5IVy4yzmoQ99BF4EHmvyYiXEtGuNbKR49cuzsdC96sKodpCu3uYqyWK
OQnzTOn2NVnykUeIMdLnPRSayoYxrtSy3kuSKTPSQ72484fAvpzYPbD2Q7uIW6Z/
sl4L6iGiU7MKLljaY0UcEweG68BFF5wHK2Pf80+SVFdDWNI7KlLZSEdZ3hi1+Es2
vpHEapKYLviQplGSNJnSC6ztryp17+jag2ZTU6ZpQnAW7M84fqdyHFAj5rKR+iC7
sqfE08NzdccKY3DnkUMEhuVGMcvEzXloKywWhkuCP9MOGlPGVn1xPkkiSw2AWBOJ
UJxFwsuuc5WmPXnc+YCREXFc0Do/w0YiHcu8TWvBWANSv1fiefN3jUafgjPfXX+O
xtE6CaNHnKuavZWtPg6ehM+0gU2QBx5dtREkahcy8gtVtirafzOTPPZihi/Mm56K
4NG+tEDnBwPnCXHE0EhtAr4qZpPNsc8R78faVns6AGnWkoSHaDPQ54YmoTaPfBzu
8udRJCEuqogHxLH0x03DYa3iKmQU72JDip7weAe1n4Jk5CFmlxVt2n8fP7FH3cfm
wX8ukOA9hNTSe/UrHB2v1KSqU8QhK6BWCfHOC/GwtUqHEc/uGhP405sodC18JDEh
lVwNAo/Hd6DR9MofArT9LOxoh6j9CNG/YBfllkqw05/O7RLj10E/SKv3eM0yai9/
xznRuJ+g4w0OZWlyeXchzUTAJqOxCmPAZxPFvUB52PvkszYK+tJyXG/v63orwoWa
rqDfheC7FpuvKRCpaHI9IpUQ0F3eL6GP/fmgKi/rfbIyqXeHj90Zn3GXz/8d4D7S
5rBDHPz/rDdSTNsMgwu6upYP98eL6fQWPlhfrZL/tWE3EP9ppNax+6PdXzxsRvEN
aT9OWCmr9DJrUkiGNeiTg6qyj01y5udj1XyIy6YskJnP6u6uiiTEPMYoNi2rjIDE
Pdvh6zmItn+PQFYnGn+cGGDAdBwSfGZJ8GzCMh3MW0bQs896KlGfa8Du4x/R1cvn
SBN75Cm5LAOGKqjyZ9vO/iWlnCpLczEpPgLmR+LFjUbUY6t0ryeJ4jmST5bZbMNq
LWW1Mi8CZR8wv5y30tqk0y6TD/gZRLPZ360ZAxzMW5fOabNODbSjHun86AcSeRTB
SBf7AHyz8HH7LjwEHjelggrFKj9wVAZAMjFPKr6zQz6YdQl/iu7jWm/fEvjvruxk
fSv3k/BQPoN2NQoFmUMGSnUgxvkGaAml+4BvhVNIQR3iXcDXRyDL3k7kONUf+wY3
gCygGlNBDtn1snmtTdYnVCHBfSR26tXBFtr8MmzZGb3UumSxPfTT/AECSdeWkZMN
QwDwDJZuCZcP0tw6VsuVmZ2iVFvaS0UMTy5HLDYmxn6wshQRwLeVAAqKRuqNJD07
G1tTGXohqW0iDgncmnNinlhV391Q+EvTRts3ZAbf96fHznfZ20B/dOmW+kHzq88T
x/P2m4jRirn7lMi4TJJJ4m5ZwhT46UskSeSLIRmXy19R4JJ/8yzc0r4XPlqhRaHf
4dofGzqi/eofrIRAB8sUPTmo8h9EawvwwxPd6BnJttz58yRdfs3SMyMkrX7IcOZi
zzKASgG3s+7YZOQjCvj/NvllOEtyCz1+Clx3E4LRBvlvrJP2k79RFvvSPkdH3rJG
te5BXRRnEo9JzM6Zsdaoq1eaurk9aH+I3IIVKm+ALiN/XIqXqo0R1x19dqxjQHDa
dnUOY2yjwE/VxuGdx0wszUnw3G+f6RTtlxOpkiyFhXi1wgOov6OojWgoUMGKnPzY
w3z3pumJ8uZy65Rmt9DcZkhUeR4DTymFoyLm+LPFxWHhBO9a7QApWYWwqwXX5eQM
Ye4fekQ3A2g5FYeZrKHM2yZdF1sU1dzqds8B0lBe7Ku7s+jzUaqIvTYaB4vWOXI8
g+Stv5rdOiUCsOM928IHKcqIygNBVsuU9s+DCZchj5knG80F8WZKqTLWTIdWtc4Q
12l2MjMwP9litUG39Bp0CyHQACPkMiRwlh1qAk52jshZ3d7NQ5YNFNDclG2i79Qp
TxRAuB2m/H+AaqvgSrj3HcuTDFHQhXCCubPeHyiBA5KRZfhfCQ9YFh+1y6WiyC0C
+rbUiuUe5GtRWeLdeYIbq4hfXpuaOYuJ0AcKljd9zDPs2Hp8KnEGMGq2oLh+Juou
C+RjQCdm24gkRpvO19HojmjOdbFlpm/QQoViprxvNmFyRX8QE0yxf2Xjr6bzHK7b
OQr5/OlWigPFN9liko4tD8jBiHLQT/oFrOhMmFK3Jq0aLW3GDCVVz4l85ZAjpu4n
kRoZ9c3dSyiZwKvldhOW+LejKMpNxd3gXiuDVPfQu7eCUrUAZzBzn7ZvroB2kzej
2jm9I5TY0XBkq8zv3ldHC/pPnuIrxLtLv5tR6qAFS21/5kDLGNYpmZPFIdyCzpSn
+9hrfoxIWek46YZKS4M2wkJc90lyGg5W0CtpFKdLrAArHD/WAT4c/wa4ZD1OZloo
okg5bG1Yn9bct5gcSZfMx6iNSAaju3fvb2P9h0YVvJVi4wA/BSK6pTZEB8615ik/
uz/znQakY6VZ1JnzOa/OUb5LBuN+ljZH1GeVXgDQHLZYReQNAGOAZxELRIE6wLyN
ccFTNGosGCN6jFF2KyRfuEQ1kl5GSlIt+9WOmQhI0VPTaZCaCnyFgwL584DUZUvp
WiHQJjRxUUlqifwxGhBhe5iXddEDaLhDouZshaF4uiCpA20UL3xVRqGh7q6JC5kS
3prw0zfCJLH3eEOPBoIE0cxgB8PYiBJg1DUQ+jIXGVGy8GUdDvyFqFZ/0k9ghLk6
ZLyna/tlsVAt55mhoECX4bSY8+C77xrNWNOICnksg+ehi39xj56WdU9hoDFSHAeJ
MPJTvgqKmhYiF9/uQgA3CVeNb0j+5CLAaEMiYtW4mvDSzw0DIvjNM917kO/YaqPS
cGC2i5UhMzRNPPqLS0CSBmSeJawE9zaxCk0mYddir/MGfEn84+vcQUCGmRt4EG9+
cJI+p2Kp06qCIRgbW5fbbXHOvY4yJRS3VxjuLnwu1w8PBxvkhhdQ7HlogOZx6KEo
iHKDR+DnWOj6mh2l78T57bBqJHChEVH58wTg1By5iEv3ekgbU257+stkpGsxpqbE
KDkpd5PB/tEINDw1zQDMSAwgwIH31rk2qY462A+rj5wQGyvaen+Y80nFtrbH9223
jsLa4h0OSpE01977AUWfv4T347yRuwx/5QM7L+WvCHwlFTecX2x5j8nhXiNIl7JE
1RAkRNEtkX5wFzxmmbBtnPQ8yZH6CYG4tpCNtqBU5Su6P6532cZIEfDm2+7eoTT6
hPaEthuhhGiA1yqvImcoAax6httzdYLPFGCXHy27FayDFgFnIOWLUSnhBA06Kk5l
6wcRl5SYExyOhwg+W25JnfB0Monjltd1/fUj5Y6ij46le5WmBgtec7yEzCqZdNoz
jKd7pTd8S7uKaU3dL/FS62Mx9hmFReTHELrPMu8E1/Ab+uvQSvoiU3T5cJPhvl8P
DsKUbdJiz7hWRXMalYJEBAkqnihjeFW+UtBLZwB8TSIYMufQ8B6KdoA2g/WbjGqm
2ZXMIedwmxVUx9U/oALvHENs6Wmvqre8db/BuKYcJYAF5sQuT2pgrTEwELAz3bfZ
6aCfwPfZwd/vT+6QMH6RfCZV6QFJwJl88VcCb8Lleryd1mSKaUGU6mlY6MPlNNJz
Aw4I+LTKIO+hiFVPtxfIHXS9qWIbDXv5KXWizQvPQSITblrfgXc7WHb2MLf+cSQO
RerG05hw9+HXQUrAALyV/Ayqw6PLjXbpXKZveQ4rs9ctSZdCX93o+GgVJNMAA59v
l/QakafwNH+POMWhMm5y81zD8KsHRSS+b9ImA8gn1CBkBIu9swphHMSk6hemtn8O
udje0eHHpF5jqjyS8CcDlXNETwJh6d38ZWhpkY5vbZRVBmnamfLrSChwpvVFvCrw
b+ePzmXEnzyxQVNCJoHvxVxkxLgj7chC/eWPZCsRAeNXn/91JfhH0Qhy9V45BUsO
rp3xZS4w8vaV+0DTIUkDV1B8ZiMoayEAXKffgh2FHk1aCyRbsycKkhW5FO1jDjCk
rfsNTxFbfP2u1mBgbJHZqPxbj0emJCsDO1DhXvZtawIsHehTL1abXrL9/uhZ6AYg
KAerRGMRkX+DU//2zqBTuZlCKMbqC0FF6V9RGeJfm5i0Xv6xu1DG4oujqIpecOfV
GNMgVeRUDkVgMFVVIE9WxYctiRhdckuPGvOXtht2QVq1YtbZda8evAxOUNJrpHaz
5ZuEdR/QdsqVYAO6yOdW0NZivry1JVGKYbp6GZwTkNgl8uv2MqZg9KriDYbq6cLr
0tXKv4mNbM8p0ZTnwscifWT8pAVJEpYSQORbjnhE9g8ykTOhhFxmxpbEfR4AMF0o
jcH5MZ5KuqBXKLoxlaMQRrR2whBS6MjxxTp5GpkmQdbVBcEk5pSL+Oe8ic3DuhCt
wL0RrkBC0WyIEPCUp5BnRE/tJZABDOw60IE3VqeYzpocgsDZBIrRBKBSMjY7T6dF
T/YYXz0wUETTsDhJyZzDQ3FHArdCXtmIyeVr73Mt0ACHRE6Go/auMcEWzLxeMWgU
1cNww0hHtGhkjHI95bbbWJi1lCBL48CaQ17+psHiOekE1PEEwltd/bENn9PqDWaW
krm98UKTJhVEXpbyfnh7lcXKxu3aXATO4WjqCaw3UZI9mioe3cTHefYiLPOJfjrG
v+kJxTFOB/XMqnIYRA5M1Ns8FK9aXeqdM0rb0p7g3/NXFJW6O7/Czeoyc/2l/eqP
09/8sveOVMhgoEnkQnHmOnKrpUrB8nHdCm6J+i8WvdHQXq8SrGAO5iK1aKozy41R
HQ5hQT/ZY0SQKJutfs46pUdDbpUKLXpvuk0Zbn0LiG0i88OGN6eeqs5+WXxRZh+1
8zhYmnromKjQh4KzORoCwOvSnxjiXj7z6GQ+WMk4Gb21luYXhLpLJlhp8fPPhtIu
dsLuUgwfX5PdFZHGEyOAHY75xi8B2vTYcNRjfLsO925BseQoXdm58S8gdHo+jAnh
G4mA2LVKQoa+MY2bqo474sr8ncKweUQjP34F1B82haIMyh4VxKSVfX8cEtdgeI0/
09TBILRYLdMAyivaGVUgirrg1tS3eTiyI2rgRRCySkgBhDbOap3mt27hMpE6BUkb
WLD/PRxWSTt7KztXSTdGA9Fw/UP8lonIZUlkVyVyeJAXqpnlabudqk05qZeqnUW7
p+wrjGFn+qxMrEwgKbWM3w7vC6mvvhn+Ww/4wHp7udHFtZbXR55rP+utpuaSc9L2
UMi7BO2kYyqO0DQrsacwv9TlqwXh4717wRCaZg0vXZw+Z9Vpdu4CDJj4Xh60/fzZ
c71ZXpsL3lPm0o1HyUIMKGO6qffu2rIVnsRib0WJ9WpdcmwB2OvOucXLGfAvZwcX
R7nHM5mw7pXn5OEc+sca90eId9rRNZD4QYcdBHDgPQ7usq6AaPwLzY+dlnvDFXXF
yOlfk116Dc4AtNLCTwJ9oNcxusxkKoY1ib/rA5oEdhiC/I74j7flIwbJO25s2Dx6
tufAabEaio5UZNwsB8VubDsC6+piKhbhq3OxHJRklAbiwrxJlonc06JsUGHuL6wC
4N2NZUIU171YwMncWcXeqOzXeJDpwQpLDhyocbRjd8dWL1UbcfLImvDaEzTqQdut
IBAU+2JO6UqxMkQoIkM4P0G/X4HUrKZdSEgvE+LSSvo8w4vyDv8Ve6O9nlypMr/c
c8hcjlTCdGiy5VGR0xrmwxxwJxpDKEh8O1YVOcf+qK5P2cbSVGp54N4jkaes51Sa
q9hBPJiAW3gOhhe0RbE5cGtnKvaa2B2QYI2WPIDyZeM/vYNvS5bbj61IOmNTlUcG
P5b1haqwDiP5LMOYl2IdXbwwAp741FTCChT9j5QESzAhuDe59KmKyHlhigXCMMPm
pDmOzreosJ7+8QYjLFmceSZf8PyZmVzSZnIEsYg+n0xVsiIB7+lobKGWEbIKloGx
5ma8/n2BTgW2KYMv/YNgB1YLsu4ljwevefY9+Pt4Q9VmqGl/KPOCbsIQzZolrNWa
TXc9UsSILO965X18GmDDCLtBGAmd43tcAZES/tvmZQqT/RgYJm5LvoQSOMq8Efj7
HskR5Ocg+9rzz/RBXWwStyxKVBJ7mAbleW84IeS49FjZ1PS+ny5Y/XYKF05yJgVB
vHVqsVm+UY3d4Dl2DGyV5TFsZ6rjbCt+5J4YJQb+yZc0D5fLnOchDWmU3TF6jpNz
gWmF79NP/GmoRCjaaQ5JYAnIlnh3idM1oqvExa923RKaIwI21egnUxb8ngFc02It
zv9nct0h5k9SPlj/Vq+3i9fNH/aIE5an/JyyNF+LIG7d492zwMpFfzu/ZfEMACDj
VxEpQx7kbyrJRd8D9kEH0JXIG/d1nEdqSIT4gZvMj16EdSyRKPoTxg4c1QiqV87m
PlY9ORuSZ93hQZpRCJu4PauNnK7vS0zCa+PVv/cSG0bOzeEme1GzpuPK2vzrr4pa
nGDytD0MaMM1wlcW5a1erwAn+IWy+xDv1kZjGuDEOc4f9YCNZvZfKu70UcEyBcRo
OEdObjDc4cuM+Q3FEB5bejiMAcrkEMk9uIB0BgraJ1HsH707S7XhZidkSVWQy/BB
YNlnTXNYheEJCr7gtWErclUSn4d/R/p3y7gUHUUx3LijBd4H/oyZLfTlR8afb/Lt
YZhb0SUMmuAUN8dezlQcoUhLgWtDUaE5uVpHc+nxzIFAcChC2U3ItRyc0AJC4dbs
EoVeETySdgBw5QMAf4WYVX9Erg1pG4PImUqp4jAOzHFyACmp36sknQgt7ALr2Kgi
W/POXL0Kt0V0HZAp6fj801GRBWqiynaZDQTZCTB/HinwvGevwlw3eRqiUmWqmwVW
gbcksus/KB1hbD0pAf5wC77K3Y/vcCLgL5uoSEokzZc23DiFDlIkXgwqdIqK8CQZ
nvdacKJJbTuY3sVdhX2uiZBPfLj6qlcGBtVT6XU/R9LRAqzsVTfwv8MIiZtChaRa
sHY3zHay2XqdJu2EsB1J2dcPKboQ1BIva9IA8ak8gzdoazy097CdkVlFg0u66bDP
LpRVk9g6hrGJsPPzIskaw+wS7GJna5RrwW+1OIrhZ/OsY2mHVZK4IyFzR1OjdOrM
4ske8hKDZW4I+XrZn/Pr38Lx4c/9n8BNwOk49BKGcZjlGW1LKedW5N40yOM3GKdH
C/NMDT4kDKce5O8+u9tFFo3gxAUDha+XlXTDn0lQMHCLE35csTD/NV65lm/5Axpb
HsfRfAxsJjkihxBNusSdd8TjB6mu+zgw/wMRVr82Aak1oEwv6hFCfZS2KCFUD+MQ
SzMvJFqMHKlT84toSAG36F2D8GpX2kvbELgzr6PmqvHU7YEgxBGGJEMb8hhRQzSq
EUmy8Z55Ij1BMaBZlvewL1haWGVaRdkt1zxvwtGDIn7uQTbEy4uHsb75imYbRjFc
frLaU/IFRnKOisZo6FEobBeY6kDowOW9cYBs8jlCqlYKXT0yQ7cpEG8AIHU79YCd
Ks5uGXshMlXGLIvZ00dGMs+dz1oYny6+7E5JJil12HpzgHqqwTsPWoQ6PblKv15X
2YwCJcOPHi4aJDVkJxO0OdE2/rRhE8a7CiIwUhxYTRZkHRMgxLy1FiOh/2COG6pq
DnX+xCA/w8++YbykwgsymDE48KhbjR48VZSBvTLPtHxWXWK0qkQN5LnjXVSRW0rT
L3uIu+XD/NOph7//KH5HFg2PRGGvXyy98HYDfVr4Aw2Cq2HJJyZwPW0adjv914xd
jY/r0E37J5h06llQgHPmki4S0dpLmEQH5YmkQTpgAZUxzxPML89LFuLwih7GEkDZ
eMb1TB/W0msbQfE8A6JBus8DqdLMo1uCohWnWvIFX7KB0UV4Q+A2erc7Mn12kZHF
NbETwpJIT/FYUFTTzkV5ku6B9dQ1Icueis/GYLvemV/vJHz9a/mCsO37lReKDVO3
PUSqMZqD9mUgYem1RbyDLzvovGxzCvmanBR4nP7c5QJY8DUPeedO8Q4/9lxvAref
OHv6rloMg7Opd//zq8V8mLzLj6YQCwat08YkSO1/ljsxuy3/IZI3g7acdUvGJqxp
YNnYSCfBYXnxF03Apwbm31K5pmH5GrFQGcL5/c54SAOpAMK+ColoFYFUQ5HX2WLw
sEuze3rRi3HRp8Xk7UlYf3dcwBU+eOkNGCYly0MNtg/1h8VrPz12m0uvbSWt2Qip
/Fvv5dwu+EGfAuY5qjobPYDAy18tEROP66exUoR0mP7BNDCK1N0APNmGi2l62rDi
tMY4sFq6wom5bx0mjSR95Rg7EGT8wkkK0Lgawq8Vuhs2PS+cpkX471rgPdGZ6vIp
7im0dJNmodGiZ3Yw+nFToIEjYNHkgXcWQSmxPI7HKifyhceEaYevOmmOdj70C81+
C+NlW4xbHugFmcgnUuwQrib5kMvKGk6lEtYfXKg6edvQCU2BEXDnkpZLR8F+AVGs
rlXHSr7j5cpqyqBGEcnGGDuvz7TEVVwMQvHk1FVFBJseDrNlOF89BlT/l3iLGCrw
Vq/DzUoR7lIA/c/Iht2CXSMsgBiPgvvNAhpAv6QJK87kloAMQkbITyG6MGLcvfZS
e0aFX/WUYI+5Ok0I5Fa6HII0z/liITO6R8wLGaKoCyv76ANAv42YdHdXC7A+E5Wd
4IkBXrxwvIVUZAaQlEWSGGqYoFEs+Ylvf+X2xFuM8NFzcqrho/mQgj3wA1MwBTyF
ZeQmqTXosB+u73QyZHgU76baiBkXnHE7VxX4ZiVO8nf/rzF9D0O+z0kvEClFQBdy
xJXcWjDoqjUuJbk6oErVKazfK5C2gG+QPeCYNYaoL1nMykf2MDL7QQwG3FutjZJF
hU5ygvyEzKHYVNtrvTGDi5bA+DTF/gpow58f0lKoOUixPgLAfOGK11hf9ttgvtDG
qnp9SBfm77l4/4VqP7cOqnqBpjl93YWTK3jR2D/EnxJbfAyWUt1+4Vzqih1i36T5
xe+8Icb0YDH5KGye5bIkaoUBafwklliNe4sNWtiqe6hb61x5vyjwaL+fd1IgeaFq
2n/QJB5hpxVpLI2SXZW4Xz1RvQqdI2PX84Zd+IG1M5DsIdL88evR3kwBBZg1qZzA
xaVVBB1hTLNGMERWHdXkAYXWaH1rKOWQjgNN3/qQBo1qY9lP1TjY3y1iIeJI6D9U
1ppPM3ki6inKjaL8bEQJ99s/Olp28D3Igtw7rh8SUm+PcUX4rho05sdtB1JcDk/E
G+KWJSf3cZDCpkYpx25YyO7VcEx52QCaASbIeq6tMVKnb3cMHDzfld3PK9ywuTRm
v+QdtYvLdRmwQxomWMgCLePs2O/4sWHI2sRnRbFx3ZuEA0ILgb5gjE0PMyEwTzQv
mH5TTXt3fcFVE3yNRYyP1NsCiPapI7WajpCyBiT13dSFQUjtJU1w2F+0njDpnkcr
Nqjgny9kCgEt1QO7jSQychhOEEloelgYOZrmn+eLnd4sJayq3FUuXbzOQF/n7G/+
o0ZNQ857YaGHXtrFBWYicRBD4noCCFyqWwvzE3GPULPcE+hylU35Y6t1lZp1kgGM
oy2aKxHUrosY2LlLzh8QnK6SCEGtz/YrjIfjHv3cWuqkbLpNhdTgFsHCQeUa5mww
HZ7rBSNXc6MPv2Bg033iM1KkmJ0MRY9AqSt4wh/n9HGvoQucb6L+F7FejaUwr33H
IuHRrkQrS7+pgODonUHHC/+vgK22+TmPLQ2d8EatBI5a/lZG2G+rGQAbYwGVQiQ4
K7I57hTD0tyISXnJkF5Pf9c3UKYQDNhomwSj+IVHeXTGco0tod4zwQxujwTlfLMu
1+q3EdK/JPr2oUQ7c60swQq4+BA6GIk20/q+YbmuL78DY0rsxxyWiidbybku8GIe
MIVPROF6d+ZDJFQ0iKxJlXNBoWpu88tQ7IumhIMphqkdmSM2I48MoKUWcXJ10rCy
KQgFp1HpT7IyUP8QQ0vY+XI9rFzMzGiMOLRX8mPpnblCU12iJ2RW1poPBSg3b59G
rMZr34lVH0evUPpYnmjdridz8LpiPRiBd+DR8k0pz+sOjGFwnC8ZEhtE2523KUkl
OYri5fKoazPBzECFcBmnBxHO+iLG/pGLX3h8mDf9D4aL3Tp2x+Kzh69KmIxn2gFY
XKrY98HgSFo5Odl3p6CthpT+Wmo5eGUvexlqfAt8yiiPK6/U8jc71bPk48PYN79o
bDxNl6/W/w7sx7B9odgyRuLFOybjZbGM5HGhBv5AelKhoJelA0p0h9Et9ap8UQWF
okpysOYJw6CER1qC7H7Ovcq0FqmRyAmpKw/1k4gwktv9ZAVpJDKzDraE7QLgaY0S
h1i5KMV6irxgOWLOBR/FohzFOnc5GjBFHZZR6Y7vOLX/Rsfcf4h9HzAmTCMdBuXp
TESZgC9GblfnVGJkavIg2IOgom81O9DxTBAyM8JLZHSq2yVk/Z7QwKWe9ndevUxW
no71CXE7bvsgs6Mom2NjO3vZKQnp+qjWlSqdF1eiWScbjKEXEskE61O2JR82Kr+3
FjY2+CY/vOykKbt9InDYAfsHRM7NiwL7Vq792OuiAAuo41hjqzfy1tm3Nd88CU5c
bfxzW5IMptTPAS9S/fSCF6pEQOkmmDutUYs/v2AsVILA+c7zYjE9QN5OZTUbtgrS
+d3UhVCL2PnQ/KbA1FmxGkoHpqowXLLrnmI2cvxbBvICDBzipf/XFPTmQEBboxxL
QPpu2WqbRw74tLqJ4UOmGUQeyKI84TvkAbrHOBbbxIxcDg9z1o3BPAdpzaVwWyAy
kytYMKqPUTapul72iNeDUHX9H/J4h8bvUQLTG2mecb8JJM32pxa9s2aENO7a2Ui+
juI0fP/09ykZQAYD6oJrlRRl29v/mG3hroI58JdWqnx/5o/nf+XaR9GITqV/fHJK
hqtWf9cQpLd5o9ptwBZIvhL4mtJRf08CtZ/Zx9ELT0IdwU+drUjC/aytlTstrafE
r0PiXI5z6CDuKvAzQQRL41HITyrYeEZYbaHFrbQhm768W4Guzw7rbiln8zcjwS2s
36AyjgrGG4nulAWBqpczQSIhkZFJUS93kYP+AwWrcVcVEaZ2XK5aw3NrTmd8M4hy
ROwbIFQc+LOwAyp5+TqrUAU+L7oc2sBKfUzWP8NK4tIto/mAfMw7ehMdY6XM0VjB
UKiPrdaQ1iZQbtJIMmBYpiLZhxWhTGqnuYTHfBiZ3exsQWadKZy04zAILkaeSFtt
BGuDOV3YvieQQcvneVRcng+w1fpHS2+KXDwVuEdIAySB2OHGv1ZxVY55QtnBmPko
pLZLjkDQ/KwpqIwB4AoIQp4vT8i7YA0WaxnceAUZaiN8nTqGa/AkX623vMOTkREm
mKXCzcvcgt4aQgZzDiYaoj5xQacii8Fjqkn8U0BuUBXB+rohfPxhGOl8AskUKH+6
SEYWrL/3AO9LtEcEL3NIGwJ6dyQ2XgSQj7Gi3GfK8z/xeKv/wXIZsGgIJVLLfv9+
KUL9Yb9FBhKfUL1LWV0M7IoHKvBQiXalEILE346S4QmsQrF3OF5mWOTQO8VMPRAg
TKasqKCm3rko9fbwbmyzuWn+LHgdEk/SQUjxfsSMA7jc8uWX+JcZW8Q+yTMUxYhP
fryjza3f13Q1NWwVpWses3skPJidFXUub07IOhFk8/I4D1WHNs8QFkrb4RKgsee4
5l0HYA+zarZgvnM9eUvVT0DghnnhYfsYdYoLA5ej1GQwz6UmuIjJ3xrDygJh9mtW
M4M2YN35TdYfEoc4MrrjW+I6NifIU6E+9/qIRpznZ4xhbtVUj3x0B9K6sWi67iIG
E07Y7IP7FzZ7cGIWIdRj7/T6oxkpz4P+s0wZs0cax6YlqBCfW4UlHwW3m9Y2WTkb
d03fh5dRsG18ft4aZ594Vnq/zmj4hl2pwWRdBS8iIqcf1iMd70c2RTylV3yUI+yr
jtKXo+VhDtg1sYDGgJWqcS3Nck85p9nV/1e/TMfAypVhTZ8Cb2wGOadagW/dNcXm
AZyjq+fDUdw1uWmlAYpImeKmECZbmnGcSqnm30A61OVKOXHDhup1y5l1AmfPggSx
GVnPCxQ2/HttvKn8lCWSHUc37qXelktGyQvNrA6xOpf+X9ECOMlLWXrdsCieAdBz
+YRfzLMD5kE1X/6q+yPAlODvp/U/M3u9b+rlGGmm2pvYsdPyRK5UMaaH9eX5m5VZ
x2y9TRZzxqjVMRGLzbj6Vt1k2uhw4s1NNEu9zl/LSrNBry2nH5vuXIdYlZn0orHK
edeRHkb8KwF7PinyColoigpTJ4puPjnVSz0HfQlsRmOK1YGq9B21jgpB+lCJAvTE
P6B6HWqlxfFmkGPcloSJLuoJDftci39qxTe7Ic+nkLcuC8nPkb0nF6bBIxCcrdfb
9PN84jEaf4oG8mxdV8/hyiijxkFWIg1ZyeYK4MW56baqF/aMB04F3XKbrRlt0k3s
h6VN9Y7HraDZ0WTVsIPmu2T9dZGWOhly9GORtGOll3wDq/MaZIDB6K6RdWOnzc9B
PLnPDGjkRYeTfLRXZCtEMXfdriRG/P+D/lwPfbUaDf/0/iAmV0thggYWfAWUiLhz
fZlkSAALWlCyLBpilWn2jeWgFXHxKHXoV7J+ONbyIqsXV/51NvmnOXqxfd0fuRk4
LgEw5bboYex/a6RUoy0DT/QZJrZXhE9g4fccAI0Qemv6/HmMcWGjgL0Ee7Xog0Ag
8kN+hy/RT1H2jYO56GnXX9dTAgq0CJviKaLDBzdo2qIaUwRXpR6KZxFa6j4+b29d
AyiyNXMO0qJrJyVIEhlGoWRwYQ/7gdPv0X/+7GwRLx24CZDFjfKaNHwPhr1j8Iwf
tcKCxgE5xE5rBtWLfZ4+o8t5fbtL0pkVUT6wGz2nWdX6e8XnGwAws0ZTbAOwBwqg
D1ADEqi8paDYNvDrOBud9hmfO10PzSe0f4tS00vDjcZBbKAJLka9gTKq+b1IUo3a
TSgBffp5ZW1OIsbS+xCoGnPB7fMV7KhJG0uBrYsC307XeHroLG4bE5slkVCP0vuK
s6PmckPO2OFVGmyhLqR0W53ltFlM6gW2a3LIlBMha/VQ7iEYrIfKckoouqziQnfe
UCTHK/Je0HDaJNsqj6kJmAVOGx9tjQ4RcUGcseqPt4geXmwAwrji5zTlKH9Y+iXS
/nhDoWJwbVfTQKE/3nBRl+Ja39V53s3m1bbiKemqPIHSh+5/z5vFVT4M0ft5d6N1
qPSSDYmimRkdoETM6q9val6kCRO9TOavnPHkKQlONHlunlCPL8EMFIPjBJWcD4a3
MIsVO53eojtcxLikJtQg9iC4j0jT/EXoN78ZTtxm6jYschVz0AkVnIXajSjcOKx5
ffSu7+rJlUJCsTYluwGEGksC9XAon/6ncWwCrEtp2s4QDnayPM/wHufeoGlFCFnP
cRTpgU1PGuKPza22Myu/FEmU17Ne7RbzD/nDuRI7wu5tp4+GPgVWdCLVc2HyQMjn
AeXRuUtAQ5D7N/RPXE+F2QG+szjikaYfC0VguXcse3lGr+qpSjPWNaZYG6EykkHj
88etCzBbNCf4t7grRZhKNjrbbv+Fu42gsWS/SfRhktS1+uRriNP1UrbT0jWhwUvq
uZMZrPmmDwNbaGnWOq32T1+DMpfc1cdef1S6KC7wjXx4DQehmPOCU5Oc2rsvgHnd
u91bzeLiBk9gFtSSIi5B7cQFcBv9XDV/QULluZDhgZIj2JMS9udWIJzrrwU4R8xK
AekYtF8UPtAGEhivI2KIN6949RF5QyVCOf86dbdaErA6RtG3FKha0bQs/NxaRiIw
weS6XHR1jSk8tRgwV6Gcpumq2HsiSvv+pMxyjRGDuaPYt7LAzIK/7aFi8yH3ICsw
AQIIpVFxl6iJtWqIlX62qYSjyyeCFKOAPBWAqD58vEWxVa+SBiZdz5axv6qmSrmf
E6HFs+eGDBm5hr1vHnBOI+dJONd6nAFShFxMhiK/4AvL33vxPtsmFA2LiKPG6j6Z
gDITmepuTV6MmLrJi/xeAxHC4Un2rmocTRG57lJPUc5wjE0Ep8V8kzchsRgG/NU1
y/oGHPWdNbX2lCzPVF8CQwZnYz1DBr6uFs8aS2sHeyj/oJMhesKN52b3LVvJO+T7
cY9jyM0v/jV4Eo07wEANxs2AKcaXGmVqCITwKINIwi0/3ROi0EQfghk1adHnTVwD
8P7GIceVoZieTGKUwf8zIKnEAT3DZt3kOAhWi2CuPnTH8m2r8xeb5noiuWi5cw1/
O2uZB9OAgIsr/AVg+R0CNlWacvNoL0crFgI9J0KVRJuepxkqenShkugwtRI0a0WL
ZZ/A/1lSt8sQDlptQdilxh7MCZ2V2ip6F5tIhSXbL4eHcsvkdhPuNVdVwy8mDctO
H6tRjGIjHxYOSunGFPFZNGXCCkKStBWq2pXQGuXPg8EnWrd4PcqWr4okKUUsQUr8
zJEk6kSFfXMA8AfSI6guvXv4tr+c8tF1VRopmw9Lx6U6rFnoGzDJsgzf9F0E9vlS
OlTgwocmg6zs/Ts3EOKe/R8ipR4TcNakHNaoq0m04KCac1R8bkonIFdR8IakyB9j
CyWWBkXpYgfhuN2Ao6IF8VJNhO+zqy5MboRAolWm4DsOL5E71edIeDYLzfkc9aSw
Lg7kjB/mjn37S+W4YuLyGpdmsniWdeAi5YUwvL6Vwmk+ZlQ1qEeMp/mbKcJa+TIx
/b320xdcMA8m/pQCAAjGfNzc2joMtANXEcwAkqIRcA+IjcSa3S2xecVr0fsFJVGB
jC9BjfVdqBdDj0fAQV9Pr4VxmZH8xuo8bNzRCC9R/mKvoqDXv0Uq7xbB8niLFgbP
I4RQZTqeexc+52NxidQeCEqdw3hKZiMIqb2FJQksWXy/G1sqMhKfav7vTu0875GC
VEhu7KhAjL7oU4vkAkUwjNVAKE/+UHbtXdIW8jHc3H+f2xnN6BJ6eIm4kuEPSnHm
gSLJ00pPHH+P1C0UwETXjOynAZISC4xl8L1i2FVjPV7JDmzeRPSMWe8GEVs6mAGn
heSjoeFTekH5GwbnZCuBhPnziO1yURceoIuVPepozXOlA0YTtVN06rdg8ePod7vO
+LdAP+s3LULMl0nJHujiY6e+ka+z7Achs/vIebYk4rxpuYchqHnZXiIz4q5nihvM
LbxM3TxLJ+0L6Wdld+8wYWZs+i8ViphMZwOkbyUsTbkPBtv87QLNx9tyJEpkFxBE
UOzI4gIUmxiRwePrXtUUKXeUZy7D0sdkc1dsQGAJOwiKwA9iGEKG05tizqKke5IK
yMU26iX7Fpr5TFTMb96kP5ma7wNPKVfPEbxkAOukkanq6E7t4iredM0c514SVuHc
1lbcVZ61omx8k5Of23FPOiwYIm7vRVCQtfgHQZQjtmN5xdGOab5gNK/p4vUURNhb
vSQGNAOzsLXFmxd+oqt1lN/n9tvmP9tuCwUQHYE0skInA7k4KkFq+HX6O9Emas/i
+sjbbctDIdiW16QkIJ5Tk6oKbCog5G5aciItQ0yDUUolwa+gAMqrIYOcUtCj0C7T
uWXb1zwSZAkoA7Xj222+qpk8q3Jw0RtA69w5cxR5niw2uF3GrWY5gJY7WcaRz1B5
LN9K2e324OTkhEwtZ3la1UnGhNR39x2hHlfSNFl8DIh+Of9kgaCX1FUHHAUwfo3j
RAZFrbqdsfgbOqARCiQRLwXgRFMhWkL69kk3lb2M/7HBW3AiRbYfgO5tq3Hx7ML3
RnrQP8HelbQtqJlV2cJp8MlvDCQiE6eDp0Nl18c1di68eHxPN4obQu3cTnGnW9l7
6gz7Z3FFc011AcM6mtfn1lJuJEzKIgHlmBjBYrduYgUAec/KMoVvKjK2sW4a61th
qPSHZJImKiMeLEkldmYb4+9B38sLSKmK6m9FmDIRqpUBa5wC3xae1KyKyTP52CaA
mH0FBmbAqH57beHln69XYImDuQgwNXQ8U3En31WwnxDzDG2Rnw9euY13hZfxpNxF
8XJIupPtv8AcB8Qmbc0hQbtIeuvVfBlr9dfCyVWkZVTHy6+uo+qxp8BvBE+Y5ZaO
ZfYaJNK/yEr7BtFe53lT/nJEHzulmYrREMCQBR3HOXQ0QYBJ0GNHcGFBFaoKBOWx
IYPoFh4gDG16cmdiP9ck/rkhnbqx9anGRPNInRuL/nMjnvRq8RjrJsPp/rQZWaA5
M8AfW++mvsbElyuzZRxATOA/86Drm6NGdFRs8fpMpFPg831buB8oVpoiPjiHYnv6
LCSW8elzHUtu99QE3Glp4DIL9xVsD5AkZph8YhgRAO0Eo3ZPGibK8qtEUdqsvQhI
AfKJrFOu0TYd3IN27InMV8u175eBVFwAI5d4xegZkHLAj3BcGi6jbfjmhUKyPk1c
9c1zyvYkT1c1Hps5vOBAythOFimP+1PvD+L8p0NtMMEZm6vleHLqnW9+E0XM87LG
BG4FPOZWBMxeuOGmW9KAfS2QMP1lSJwL5ABjG8m+SaiB5B6bvzudaCym4W0RB+Wq
GKrh6uDjNnMrn3bNH+F4dn1MPip1x8Cuvs26OPJgevuoTFvKypQQz3W3onPNTd0d
ZbVjCi76FaSTCkKOnqHTJ5EfCBmwMxRMY4Sg+36YW+7YKGy3g73u2kozLh9wOLaq
WhkoNUmOy/BxZywjxe/CR+fH64YNWmnkpbWnRlNM7tIKXjvHnsrAsppS5E3rpcGj
15TnBiGjAz5N346ZhOXlJZ9/WYpcu4xkfcoJTDKZLMIj44D2zZVtu9nk1x2W2irI
HiM1hXai8q1zO4VNMhlrJbV8yvf8wrGC60gvM7GUQlzslc9OOcbexc51Tw6PEIQq
lM+WzPVPSo6djzkcjNZGvLaBX6KVEIo8AZUX7KtfJBGuXxgSdRg9lNxr7J/TBzKn
8EQkatVIMeR8iwPBYRF1hiIGUou+DSH+GwlAIGXA3MkOO3Qx2mNdf7DFidKOl7PS
f7Si8WqO4KJIaoxWl+5BrbGJil92sF4qDnQTEuJjZ9Vk/rBxdMoF0yM+RvUl/Ikj
qp8L/0Axm9Eden5/84tlFM0gBQOYQaUsUhmLSGoNZWccSNiadZiI4vJ8PmgM5j8z
/KYEz5PYlZdxSSjhFw+S+eu875OgFVBouJUBizi0AVE/p33NqmWFAdxrkMFBX2hR
mrc6z+KNBB4BoPe/XX9tPwWEawrahg91zSsfXuJr9tKYLr/in4fwCFiQUw1bPyNM
/MKLhke+7ec50A1PT2lEV3Z/s/flJuqHjNi0JgqszLIxYwTIPcnZm40xyah73ijg
5Bvpzy4CTRJuq/l18Jse58yk81NrNtEt0DNyyeKwqmiayBa1J/FC7WBLGni0N4zD
osOZ321+5+oBx75POSLECCuE/PPb6bILXD8x0jOhKJMhe26inauAzxhPCKQM8ecv
syfUpzoG4SUtv9rshj+QpGzyrrrX8V5BRg+Am+rrZUgGOyPcwAfW500wUFxBjV8H
ty1gVPtZW5VK/aSC6ZCGxTYhs45gXulj4VwK1jHxwJ7EtZxF702KkWWkIfmdONY2
KNtGqt3T/dhq6KYhszs7Jo4F3JFLku53MwRFGsQkFHCrF37wuw53ihHU3JaDboCi
GA7CgKbaRCS2kh2a8EwY/CFwK683rmj0Z0Eh5CJwPjVlMxAg+Le8fLwI4y82NAPb
yHQdyv+k9/4UeTKdxjMlfy43cO7NxQhfFXV4NHkPt1pvhZasQbLYnvOHT2ejKFhI
LmXGBhnPzkeJvWyRW/Ywv3GXa9TgZBFYCmqjQKNdkcivXmpYpn+sTAaBz6G1TOHe
upSO7NEx6ui48JHQrUDs5nE3zDUKOBCcGmgB08JfgeUmLVusqB9vP+jEGE1oLfcv
5VFXkqaSRagB+A4CStx+FMuOXFIzQdzXfmmR3fEIyV4YMiYBPiJXioddMoXwQaXD
bVx6fT/TE5F512UWmDc+RM7ucZC1QnErxl+I3KOWBa6s6bFjPCAKmGMhR0txf1oM
sD+iP/7fW6vfluLIMMJkiMc2lzcM30EXTUUYoJzi8ec6O1Esdm3VtyU34hhLIW6s
ysQcpagu5jDX9NVFm/coNjW7nfjyAuoxOl+7r0LZmxzJXUURL5wI7a2BqWFG0moK
cDqy5Ts2GhJahZGRrsGnlLB0Y+Q4vB6OzFCc/PH33ePKbe5ek96zObjeceyGnq9f
ctlRcSrzALw/xXerQ/ightKaB0vB+NQZuusnA9bGtNhr+hOH+6XibiKeAqr0hjNl
GtMMZ5k6k1lLTOdec0AEiE25aDKo9q0AZPxwxPXcCHVekibAelBc+FeY548K79bk
y+UYsufk38vHyoFpZMzjhWHbtNe1AZps/JQcTwidUS2mrAFvr2Ufi4JNqlK1J7rK
rH8Pk4vyuU0PYk+CPTV9JzgAVMaX4d/640nTDFLl3X3TgJQxCjAWOVIP2Az3JWP/
sVOlnJPzNpo4hR3ZgLY96lGTDWv0w6eS3JwiV5F+Ui8dwJHa2F8gG7Qm2yv/7lIm
njPd2c9vtEE80aUwD03WNSXY7Gy06aFW0evwqQ/zIXMFWtuXDsDWgwZxGk4NkK3A
9QHnQDCMnCjuC7my905sxfoHVlMo4Xmoqmv6K+zlt64/HPqd3cio+A/C44fNpH+M
m3LajF0WJ3bqFVcnHsY/ovOFOboeKLFSTMxvh/i9NPn/kpRlh4rj08s/msS2cZvD
seclDEJzrpsYpIVxTxez0eeUSABuy0A3MUmZMfFgseX8fFLhxWLTgHiL+wExcfwD
ofSIVXeTlZkXrkEyb7saHBjzeLHC01jqh/92AoMlqOGg2u9AW3HJni7fysexhp4c
OFZWTbwr0apHv47AiOuaRGuj/sTuFZj9r+HVragEvU7LlshdNHEeWRnLVtJmKjkQ
Zx+n9bm62NDx6388maH7JKWqXUyYhIkcPQmwIrZ1ldq1UVBR+Vtl+oodN5DSODcL
YfVB9uFzXp6SQduK6DfIYdXNrCCPRsjpNzE7r+uNMsTDvsbFjVAbu4x4JX2Snjw0
Dt9CCRcPpVgfneS+FKP1a5SDxU+mBzFRMoCMjoajxTkISYNNv60h9yZSnjpFYD+v
s6PLem8RUcXqd2Y0zWl1SB/51jaJI7eszUKEXxGTfxhikShA9PPTW1vA1WHno9B6
zJi0r6BjHsBeZg2fB0fMAtgzXUqe6sX4Csl6TUgXan/J6TMjcVXJHza7yiLVhUZr
aLcdN2oaHin2FcZVdDd42rpHCpaDuiyc0zaPI/YRbhwcQGMJwqFX6VzssbPGQ6yj
CB+OlsXJYyw0LtFF4ajAZBDLaqbmbf02yCD5DeBkvQGR42e44vk66cyOqjnfyTuB
6g8dv9NIstgXJvqQ1QTJvwSVULtJVbgg+2PvQZx/YjMwFXWPEfRfFIvvSXrAdM6U
UHRqdSlCkq7B1tsvzfyQIMnUOCAFVo4LkfXEGXJuMTfewqGXZQsvN9xqZ8ANdFnr
oYZrxymaB5uhMoypdcVhh36hukpUNx1bs5+cTZnLr8EIkLt30lNfNOE21kMWn5FR
3nESyOcrDjkj9kjPkCw87IcUUh9ogUtlYtLNE2EDEiIRN4UBhcIYi7e3pxU9v1g2
xiVMtebkN23wqaJlnarxkjeKCldyoLCbdMS/leCL3oVIjy5Xn+3gOLLOUxyeLH7K
JEquGs5V8peXImTf5Q6n7ii9gDcGBNtuWHCQOLmHQ1zZoyKYnNAx2AjNxlgHm1vK
L5UOlSNfER9qNZWGDLpktuIiDNx0hiz+XWkplh1WU5v3DPvbfqfPsfTsDscv2H/7
kjd23WFDSP0qQgon1vcQTb/aUPjhq5x6++jCIu8aKcc4PE6H/svct1Fi/9fF3SVr
ywoy7Xjlhuk/2TmXeCS6D92Bt57zpMOxEtqHI59wni007JO5uWsvEgogeWpsjs2n
TYRzcZII1KMzLjuoJKXIxDV2qz2/ioeQCkyxNbBis2Rwoky6J7g1Mn6OaRJGD9Ka
fbtFI3mGMn28kMGPP+wWe7Lq4GVrGclJIG0FArWK5vXJ/dPpDWbzAs/7mkduu6Xf
eHjtcVvkqx79Ha9jI3jqY7sdGl1lhbAuRLjJKkJtOqG4C/d191WIYeEJeGmwUY5I
dO4IMACWLQtip+5vov0VhQS43nHByDt3kzs5DGAEEKx0uFNEe6u+0AK2t1JWUAyL
KVGgx8MJOa8bmpADM/1hjNy5w2M8TSUZfbXdh0+QPHQW1UiysOTDfMrq92NcHW82
WSWybKf7c25m81sFKOe3cFBCFUyy9Ce+Por7vEP8GYwP7iZNWAHXvd4YROptUGvi
Y2f3zgduPNJSVHHYOG9170PhBwWPhR2JUhTVfyptmS8/ODJ4Lwvv2z+bA/2EY6xS
2zPBWNhj51LlUkfp7xFlMhJgfDPkxT4uupG3+mIjuZ91/wGhPVpApyCZDb/Dgay7
bCwGYGJ32nhnZl0YH1f65XSor2P4djTHDRvkGxn9odzVLAF04s/H4aZGbZ2TY4H7
Ju9zk+al4FeQScYSknScLN2InyjEQep5kqo21rd5RlSxgZA92R3cSQbBI36Md1hb
V62RWlZUSGN9qRmc2Aa+4YrKAiZPnR1dBcxsRiiVu9tB4ReqVcx35slypTbbB4pa
4fn26lSjoBqnXkIE17DCtm8Cp0j4eRPneP44bkXpD/PXuzz4A8r5OJrCriCnm5Ss
qhxBCSyWYvmAX9mgaYAqj1d8KkLRY6GGbRKHYI7pz9z3q0r+FN7YRtLd9TFYzZ18
WQ54opuKrpZUNd64MzJyfsZipwsxwdRMoK67XIqAsT5UJqWY6lzdyklW58sj50ri
bvsg1x5qXi5Qx81vFjb2tumcJQOu40hwk/Ii/HagqjDfj4hLvyjekrkFmorKHUbk
lRkK9HLMZhZrA4iYmnf0zHsIiXbxZH+y3uB5ZEQDBlxdvNuU1Or/vQWxnD1yzin1
51JMWUoAY/tOKPn0vw+DNpm0aSTb96BDsH0ZpEqmhVIbrCElyuZ8W1VaY5ivDl/R
IOWqXWEZWsOiHCPLdttL/IoT3OpCcqsqQC1X1c6aGn5MyfDABp0mD+XI8VIrgDA9
Wzkp04pshcCJBE1F0busgHEdAKHfhf07354VVOCxh9YeAC+4SAaIo6tcNyfto85i
rqVatK3d6s2UnLcjH1Ti2swXg39hl0R0tePcF0aetHs4ErZF+Egzf4txaEF7dsSr
AD3BjWP14NHg1rYfVbuosQJz1SQAwp2WDHqd4F3VAz/m6okl9hNp7Vwk5c429sr2
ygmB40Q1TpX3FZiLY4Flvcj83muDQDoceOUqviy7y8of6Sfyz10M4XTuPpPybI2n
Jipj3M9ykf4Kniio5wOPgurKeub7392gUlRO9gmhpldR6AZvDgYrzaia+5iyQD+i
jfh68JUMvPB6TS3lIFA06DUa5eWQqFlmRRuBRljRKdCPWX0+F17bUvkzPhKdgwA7
TBphhjRHmbGuxU3qDOiB28GACYnZERP2mXhjdwsWlUq0Y2rSNqeBQqdLGg/xmJk1
VzVrx3YyGwDnd7DUtIZrwPnow+PEymqA3QBoUXTx/od/bRcyBapkqk4quPqWgQx2
iWMDbHqG3bu3AMWqYdxaUtH7Bk3x/L5rzv7f/DA3RXcmtAjLG4un21L4fg+aN0B8
QVwalwk6wSbPOrDwMrpFgjNsizBGxZqQv6aA2xv2NhFPOOyQmumBGe5klMmnzoHQ
MT888/99w7d7QOeA14tHlZsWoPen2srR+8SYFTv/ROKkGCLSmlngLhdupPEbvHl9
BkWcWF+7+6zRVOyvnUVslqGJoC7TEaLvjXMEO5J+q/aW1A7dLnXg7l+fplEGrDzn
ImcemA2f3c1K/bEotUT46P1IsQaX/bKzna6qO5fVHDMUhM9Dy+VTf+KkiZXFtzdt
is+o1wh/XQr16a62ivTVlIYLbezZkqTtyzDA5cNSZkHyNebGpkS95emGFQCxtzkZ
zf7P+mB30SBacoQrKS5sXvx51KHcf3XPk+2Oi8QMsjaHA2hn6XVa5VcgFkvn+D95
fo2xcxuagNk1SAIMK264ZnqFoeE3TxCuf8WrMpQ7h6wXgBnoA1Q1QH2HsFR3kL0T
1KjqAyEOIbdaAbmAXfw5BRoAZTPePhoEh2XQkaZMh+g6USMimZPfsv2KgJUg5TFy
s38rUzDTerS3VyE8xWWuf6cxxXiyHiG9PXbly+of2jlr0twSR/7nmXe6KbdNPLCB
jDL8beoJPVVVPszuasHB/OPvziiPQ+sgZkyZe9ewqKNhG1Tg/NZB7L5UEaWJe6E8
3BIqacKZktSSeeF0C5zJzkGQTocj6gSxntaM+s5PH31KOaXKLFEMM482FCcpc8i1
OCYOwU1F7jDRxo0Afi3byJV24kgQ5cyWzgCdivrpggkY1uZOTRWtUlRVLzwOWfqG
yQ1H47BHwssZdWbwHViJBy7qiEyc+SmK1G+705sxySB4ek8ngnvViXx/D0483aeD
y4tBI6T69S9b4DcgAYap7s83qAOv8HePmGPd03tR4jfLSTGyWyyogZWBH43easZX
8Jbb8sdJL8bDeNEIBXXuSaYNQtcCX7onzQjXCafzHXNFV54zmQDsUX6AWbWJcbS1
aKvOfXl8Uoq4P3uIDOCUu7dAVrHoWK10mKDvFJ5L9ssO8ZmR9Sk58n7Y7GdzElbM
EysbsfI6PYx8tWxWIU1f2LyaEzSx1QhU5sVXhCUlTWA/SCWOjPtnSlhZJ2CmHlyG
8kQWM8V0a2JWWKulk2yPk2yT7LcYt+xp8Czkm+w3iXQemTCx3ynv0bmCc0SNk3tz
qRoN0QH6prbXrqnnzwTQYd2CFBWXVqdj+Mqjx4KgbiEmTHIP+qj/oDSFaw1ZZ/Hs
jLaClG424SWQZsJLfnC9ba0RNr2loU97tf0J1lsIF/cD1gjBUDvwN6qujHtGFzPS
l1qfeFo7F7blTMyIswRV511nOcYqes1yQqDT6ndTbWEZ/XvHKCqR1sYEl+hEm+Bf
BzR7oD/gxU+aYBdt/Gs/PpY51++oIK7AfYNEH7FjfvbbU6zTIj9+T/pEMcpQz19c
y45+sWQiJxZ57aHHE5b5Gu2AClq8EW5TWJfyM7qa9Bf2odcE9Kjc9kyQw9LitBlA
Ax6NIxqAMmMSlfWJcspyYbFxRR/FnAyQqtST0ka6TMJm0Ez1ASxEyCHFbrYpxe/d
5WrEhuosYONVdf5PBaeboumPd/MK1pFPiD7cdCz/QDJFew2Xcw0WCLKbmHDUz4nb
kqmuPSt9iiEsm6ABssp8XmjrGLl4wRVwQsdP/qtccrC4QxrWgPdun5BZEOnCRVe8
1rjmPci5p60Sm9pS5DFMd2SLLrSyXUg69aro0S5+pTiSir9i3EfUnDHXxGR6X8Aw
GzOIwCXm2YWJREVfeFCxZhTY7HM+QwgSvxnbQkT8BpEkTtW4+jC8YPjYvMqDe8mR
Y2xO2om7Er2mZJbirADQJXdi6c5hiPnS8gvIDmkLeCAdqlgw5Y49KhLBd/CDnBaT
WpIIUDLUbKKx+jTwBsbuZf4FXisuFCZJm8UDeOhIwbCZixYR4xEzvWZf9EhcxUiV
pSg4UM6hBKSrUU6LQgcc7gJprBUAz7LgekNPNQwFpG6aeUBtwuLh3OqMnvi4wiur
0hQD0S1CH9Gwjx/SxgmfUOo5DWqCz86BAo2EiCCTTgWY25h63ZI1Rsa8IKbKThHd
EgN86J/+hJycUgIGYpmUwfICieRXzOw/QFK1nYOBmhAHs3kikXPTS2tq3IguHWVf
ad7F4j+twKnlK2C8GvmGlbV6IeQHg0Ft9LAo4l3lr3qNbmOUOcT3UFYJGrJY13Aj
Ofv/yyc2vFko+z/eEKY+0xPH94ztZY8Ob2C+mhLGr5OXf9vmp85tri15HqrOH9X7
3fXyKUKZ8m0EbnyO2KX3rNbyhA4YsyNqXxrwWs3k3aDbXvtxudMwYYlb6KczrrCp
dcQlzFnjCFuD9Ju9lsyfBHgYphX0He63awd9h2+u6/IkiMagyQaKpwYHik3U142u
ysemWctwscWpG5Env6AFHWCEBLA073IReBwQUAEvOhHhcUFt75ZyyFvZQwQB+lwq
maG1gJ9kFwuhTmFugzoVVKBZo/Zzv2NtwEihSOpJ8Do1FjEgjM7ZfAiwnPiV/ENg
4zbqdR+B0FOeqW1HZjCMgQ1xAgCWCX+lEPGD9EUMeybIIOpAW21Z0D5aYabElQHP
3oCPBe9P8WHSEFes5+VC9pq415iygI4ifgBuRxLkidFv9Ch4XTvy7i01txXvV7kq
7hElwWbhxyZbxQwzloQeOcTb67GGYD4UGe38WdVAJzwaA8AMl5E6xJHkbklOb7NA
VRROtg1qfP3hFrt2kt0Ym+JOz/V//nQvqHr0rRmCBU8qLMG8oUCunJ0/tii9/JjI
QCtFK0cKGbGj6TNTRI3BtQ6r6uECrsVjvqNnNKKCYm25jhHn7k/GckaOUYBFO6jF
figWmyek9c5oCB5z+IsreMUX+mXiiEosh2eMNmAPJtP6S6U1zolIZpXCmqY8f+6j
8EV6bhHfnssNCKRHXqoTBboG2vv4H0ctLTiCzvH6rq2x2t38v2wVwTMOTTTnspO5
Qm0bFq+MSI+9CQaoVRylQ4w9GYbwpFH4PjPEJJAKQ3kUatNObEkimZoiQkJ5GCfZ
TobiRTcxmeih5bAesqUC4SmR8zCdd6GxpEA+0FMmyA7D2OPQzXTpCU457XDsezro
YweWEioJELjtEbi3YvUrGzPD+QVYNMVF785YDPyCwQnVL8Rc2kynR/OTgNbslW5u
TZMDiPoHW73WuI3mhvUVbXUkiwy3frtdqcFzyIX/TPIj/MnkOrBlbjU83FCKZPhc
vew+JlF5J+scss4MS2R6GVrTuYqhV6bwAos3qbMGkTlSshdZcoYGmRqjN/q1rlOJ
6+d3om9E6NidDd2k3hl8zhh5/doABdGWdbHsZGj3Hkoagf4jz8eZYOG2zEj+F21o
ovPkTQhK4/y4Kv7x8aqdCgK7H6NNSWOGrjuctqOFdozrflNtAZv3T8/9WhsPYh8E
Sze+zNBVB1IwETJP7b6Rhw8hgswRYatplgpA/oFxfL5beUBuiNgoU+RC4lB9/k38
7Vynhxo7R0Td1d3M5l3J/ZmfbFBsgV3nFG7SHJeGbnrVa/UoJ3AUVaHmh1GHnjjB
Y7K3w0nxcjHSNXLlrjkRLWPskQMR15iTHkgXQTftJ2diEblrxPPA9Fu8eo2/99mZ
IrYfp4IO9p7tIvFgnDGSDaoNPaIX7KwUc1ZAbgG/BPFLbCVGHgNApClmuX5+X7Z8
uL3f9RPw5GTpAa95l6efnxz7+k5fdah2I5olOgcFhelyeT+NSWCpQEB4JUX2VBpN
2HRYOgwnGRoTtZZvizIlc2PXk5l0CvwYzccIHuVCu154Yxx/GWZD68uFpDtPlAY6
E6+oADPhN6s1PzMMrdrW3tnKRl1P2NwNUuuU10nf7GHoLiAgaMSqfzUbvlHc+uor
kL4+NVHb27YgtF4KgsK3YjcZ6fB4hsFvkkVNl4W9xAKEgYtrFn+89fodt7qz1SvD
mTWjDC0e8wpwsACO7WfM86FjvF+LldpEmmpIwFFa51zURwvMnW80EOHGT2E3nk7y
2vtzgoDVXeZoDkhzL7lc6JAF1qFACil49PXzRx0lMmweCVbVExsjhJe/n4p8Cf0N
IUL8EuuTDonQOFQA0eAPWb02pZVd8kWqSEw320mz24kSSXLA0Lo1CH1dLbITedi3
ZS5qrFaIUX6VrFskwZweFnJOtautRpp53fMZxU/iHN18b1WrfSxJiyqa83stTjaF
Ei9vhajgm0lgMtDdRVxEMzZahFgGdt6Z0Tn+bDpOaFBvdFE5HmjYbzkC59gSECUb
IdnEvQkDRuoeq7kwJdrn4G4Smc3Grmp5ZaQ6S7zsfARgT3+Ic9pPutumcVFYHMLr
PGQ8UBoAQ3eTF5huqHToQwv1iOA4zxOlsSiMZnWjvuZaeLcLT3jd4naCPgN1hfmm
I4NRCriUhOqwVG+5C+GVvgv4jwKm9EZ535uj9ACnmDLh6hWGdfgN+zpn8umdnkjt
nWSqP9QeBcaT2ZX4eHrOpIa5tZhYf/mEyF7OnExoh3/m/A2koqTS8xE5+BMVF+jF
MJQMFmROEjGKvrnozHLkZjg+3TqCdjh8UtQ9bJCOhpLZo1+NRjX3/bsPoEr23qrK
n/2XyhCTlh35GytTFlJ4T5FsgBbiXeryRj4YH4Mw79W38UM5Dz9kud1844xp42y6
CsKgp0EZm6mJyaVGLCow0fpCBu6VplQU7c9WynjBq60M22dpM3Uwa7U/Yp+J+AcJ
sQlxT3a2TcOcKZmpBf4HYSt4ybmeMOWD+DAr1uUJKrcmX0Uv1pqpnNdsf3sD2nir
Fs/3stQ2gCCPlptbNonHsETABO+IBJ8d1CGjDpVZ/fHLeDvauLYbqm/yJ0/sQgkL
3PxWayOxoxVp60eR4XzVjUNP7yqF16QtLH6yeG+6J1wSHhwko+aVqPv1zbsR6yCS
vP4iicpLe6rgdOIiemeGUzRB3jvYZAGVB3zPfJC/qL2+EmmFEisOa98M/OA4R6f5
OC7ta2AKHyTAozA9QkoU3/EgaHXkC1pXiG5iK0JkBRNB01mcaLKNTk39wpTWx+Cp
kyQOWbkHxwOWk0+4y9YxJCFVhFahKa0PQ3z6INaa70CKcbiNFkJDmLipgv7jYIHI
jlHFMr5yPgpyQKhu2ZybTktkDz8omSJ9tq2Www3uqnshNu38EA0TMvSbypd73Z2d
aKf1XB85QP5fz2crU04D4svbn17yKBoPiWb3HFDpN+BagkSVVmydpENHDYpvxjIH
HbccH9AVH3bbIDLAG+pS6/s2t9GSd4PJGGVWOf7DGFEEnWQlNMoLzHV/ndDY5f5H
mYzunscyj8rtM2OLCA26TfoPMSRXwOTNh5kuQIXuQLjQGKvMN2NwJtVKk9s4pzD5
DoXPAonKCoByDb/B3gnoUMsURJWWeO1gyIhO8tQ9WJr/HeX8M8hCcKj0DH9JXDz4
PH5kAoateeVs+HbDO9xVOe+CVaIVH6FLMWgwBO4EyYmJnXMFZT3S2vKIuRJ0rbx4
DF/sAl1/xnc/u3bAVMLY7NnFyVEPJESLttFYxbzXPmWeuGwCarIUlCZQbQ5IYk65
PmYAc4xkxPIxSiBZedbw3/RfPSFl+BAj2tL4rxUA4AzgqfQJgVvE1/RkeFtly9bO
eSxXrrZIadBfK6EDPKFj6Cvufb/hmPtRkT3pdnm0Pz+3dbFnRR9ovr0wXzd0iN/I
lJdaPYZ74AXczltc7MdIlu7aWadCrokVtz34n+lL00IC5EeRMCUO8E+ealxJOp+4
o40ktKCu55t/1MGr79UzxTb7S4/vUBNBcGMkMcISnEEqf6btrfM/jhJ4f90lSTeB
z5dQFxG1yA64Gh1088EV7yiuvHk3DHQX+lSUGYvrdVm1FiJbyddsKWjrvFe5TxOQ
e3renaiE0u+RNNoAapje+2Qr02lb2GoCrjcYwBHKSxypX6lrOl33F5/JMjyVfqzO
ry0RUzy7mmLqXz6/tAipYkWI//xQBWrY8N1HoX4Lylpl01PGUcIrjwZcNybwwnms
uhNKUlNDdPt/nFOADcR6i41zyO4FTnb4jJEIRUORWnjjJnjLxQX5dh0HZ82sYg39
bffLEWYQpRtU6fXVsXMeUPSnibFINKXY6VwsEMKPS3ViWwJTwykprcvF308XewX0
DBYCXZUS75tOyGy6o1TVJqpLMsW7KJq4QKcD781Kuzk35wLf6hrmfDtwFkOstLrC
8TyVNmSb+bumYs+HOuDhIkfb0xbCqNLrZU5tZ7D1T/BoDbCGCzC9Xp1gimnwDQIC
7s7GGp2OvStaFkX2BdsHXbMwLhlEGcrBEW62eIbjNL0fdXBUAbX87EzvtWHCbA99
SW2bgz+Qyl1GqMfYHH0as+NnnzjSnRr03Wu2/EP9JS5v+MwVxf4BxD9+ZyCR9Q9k
vmtn6VkXvAAinRA9ou02O80ZHZcUadbNoUXrsWwdWvDMsfg5vLFaLF3xyefA7ad/
8mMg6tep475ZVcC+rCg/drmJhxXIFpHDfaOaQL3xIqkX7iKFNGq4+g+iVJE7jXdh
rNU64JIODje4JtjsD1/EDYQX7ofXLJ1a2RP9K2Z4R6dMbwPh99Vtnqyx4gTQHaoV
I92abLK1uxEbHp4Uhi6cOf6Bli1F37AMO0eCUc7zSissH3SHQWAeYQ0UlP+aVXdy
MVfyMtCj/v2Fx9AepysSg2yL03BPfn5AdRzLJ4PJHfosb4/ijR5uaLnEaTNmVhpM
gUwp52lmKx2clyEuO+bDRgDxRqdKLs7WegqX4J04P5KhWMJSeIWStatrVfu5BfSF
VuEPn/1sNt98PkprZ9RjxY0szd0rTmUHB+nPr0HR/TCiPrLFngURjKgSbW8KJKQt
KTInCvmwxd3CFto/hPHSklnq/xW9U0MWWEoUzev3mNAWZe1XOTFlzNNeeVmx7jKu
B+1vsLt3AUXHTBZhHIRxhRQdXcoJW5aKBobBt+g94MoOPC7gccPjiTjs6ckQ2qIG
FqDqqwijGXtraodvqjqk4XBlln2Qy9ZziPLTapqzlkMQ3MOWzwq92uEYqmECOlMb
9CxygHrj5Z9lRuM2qEJZsyusL3plwPvikykxZdrr0m+S90jhrX4qz3b8Z+FtXR+f
a9cAeyaYKrTG+XLS9Y4TkURL8xV9pjTdZP4EIEXE+Bf8gECzPcQ5e6pST24VVUNW
pzhETbV1vdAB6367vrQNaMV7gBXe/fZ4mLHIR/yUfnoCBkrLhxkmg0A2NfeeoUTJ
cwlAdwBqOypbv27pdMZGLsq5tWQjMsHX4CMzPb000xc052Eb4mmRHXeMZF09ELsD
SDF4TISQRvS+EdGcWOer5rz7JcQhdJa+cYhEAyjCMlTnDFbUqxVqI/ub5c4sLHu0
jwZxygftxELTLN+a8+XdrAWbuAOD8UPfQge2Ivx/WrqMCkLi/4izSGxCPjD30+K1
JnvJ/Q+ifMSpIbCgRT0CV/+tM+ssoIaEdmfzC+XHJ0jgIZgOTfx7F+jhN4AWy7DK
RIjk0clgyaZXpI6jpK+zZXIqps/sxS1p0i+4JhdNd4dhsjL9Lhk0Upx5VmEtyozo
TCpZoBjZVtp/LG0AShI7BP8NgGngKxiteGyiErfCIvo5SBrt5eFscH93nNScjL4J
vcVco3CclsFl/4wU9U2nA33G1yN+0Vvgoh2yK3w2ct6yUNNzABDqQvD+Nn72FQis
L1/my7FLMENzIlWzukk54xrRuJa+0vzL/m7pYC6pWfI2t42bMMbZ3VK1AMmmtCZa
0pUQE5DYDp5MG08vhdhCMJp7EEunOULquzLKmt1B54bC9LMfJtW8C3Q/47WBHiJI
q+pDQaB1Ky9pSVutOrRMllnViGnIWpLxZLZ2v440wtn2ft58yWLbI0LmgSO8TYkw
8EQP1GfRelKP8pCkKJl7U9yF83ounrahx2ov2FwPFcGe7krDi66maiDfNhmkEaOf
CI3GXWYnmInnZ6d3hb6u0byri3vA+cRVtkrMWS7PldvNs1VKzgEt9d8xCmyoVYEG
nQHcplnwHBHc8YnFijuYgDyc9fIotzeq+2ckXT9h99uhOYEuk6Va+ZUQxGPW7fxc
qEv/0V9PUCQBI1XE1+Uzv8qsas7iTrFt0yWFuneeWRZKaZvQBMz1PbnFiIum+Z6L
pKLZc/qW76/+7NLn1kfhX1RKXRbUilHIRQEsgAnvDTgPOf4NsztXpiWNyQFonLzo
D5wiYge8xbcreG3fOd4SE4timCG96fbKzM8YXgMbMUfECZvYtPuObyY3y/HNJbsz
NA50cvVGgFmkDcmEa6ra8GgQsnbLX1M3G/ATAcOuuqJy3SAxta4jneIE+7gdeEY8
P80+7pv/LVrFJMnpFwX8LgMMhYnFHVdJsCLSJ2acFgKuJonq+rW/Suy4PqdGLzQR
D89/Ec7ElhNYhgjzN5B8pENJ5C5P1THMSd+D2vnrrDRSla+e2u2ILLakPe4TNmXw
7jytgYWY6gQZmt75IGmLXiOf0q2QGMQxrIvL/BLwhsonqWqfIRFXt03lxHklZUZP
BSRSS18DdyZLeESRppBWiKZwUgaKR4OxBpaVUqbCJUAC3soe2hJp9PKWY4XPL3ad
Ljq9pg3W++Gh8+EVzHEdkqh/pFg8Iw5qsQYMKfs+cUlAi+LACv8gYXRVlgn2aYpf
8bcZWyKuUddLYugxOlRrt130C1a6XJwRoxnTnfF8LDK1P/cqWFljBwkzYmFJGdvb
wCo/SDkKgzYucxvLKd+LkmIFsUARSuKWDYJeaUgKtlV9YIQujzAhzsd+OQRmS1bd
G9DMmqYGkITs3NZkbtmTVqDayS2dpc5XNOsNVEf7K+p1rY/SKk1poFIBKZ4EdzZU
AoUe7Ebb5+ZGkLIQfK9BBsI/Q6u0MAWoS8MgP/xLbVLaqbF/FhmiVOIHhezJRYuK
kkSQ9gOpZ9k//qkZkShkwv5mqb9xwgJZuNSOXsdrMdjNKo2o+hrLoK3ax9Sc/3RB
p2MvOCHbvdqdnYDrgvpo6yhhypVXX5cRem4C4r1kcfb20Kj/xa8qcgQJDmPU2KGS
bsib2BloK6GpvvRo8xNVYAcbyEnr1InQOsWmqUM4VsdJvvSSa6FVVREQ8lRIEuJu
y5MPEWM4BwvVDb5xKTlvveK7MBN+6zwND5tdm33wmJD02DNsxM8GSc+WHXL13YgP
cJYqSUqHbJOSbFv94wwSCJnBx1gDDpvzPY+wuBj1T3bMIeL3z8mR9X5nQ0XZFyw9
bz/Fcgpm1fYmDu8tIwLMKj/Nh7WG+9pxT1d80jl893tGMx0JUW53egUmazdbTpyI
ocEwF+lN0x0FkvQXy+whIK01iTY2KiyrzYxrcPMXhCaXhbWYkvX0UAnNTPrV+Ais
cQo2/KPxFA4e5pILdQBC0jg2qZp3poCMTLeUZNRx4FRxSztX3lixy/Pt90kvEd8E
DNuJd24pNlfKsuAKE9ay8CBuDQwS0oy6ZXRfcGq6EfTmQXVrrfzqLe0p584mV8Up
23u1X0eHcU4tuZdH0NWZy+cci7n697Om3rPyv1bn/E0l1FuSL7nZdY03q2PnTjkl
X9zeI3RjpNQ/oilqPRp9V9YlQ8keQeVQ4CV2F8Clhl+HyjtYibKtvYYM+Yl65aaL
fZ2JQ2bO9AkyTcR80Ns1AC0aEuTPCRO+q/Lqt8E9PzE0PKpFpO51VGcexdlmvn/v
0YVJPg7uWPgkChdYuVo04x5z8MSBX+XQ8r4C/6r2fxXSGkXd2QapILqjmMpLmIFj
qew7GM+rnX6j2D136rDE4hi3SRXAK01rpY/+/9YdKKHK1zrqGsKHPLv4xWpzISml
Hxu8CVdFNWfFTXpjLuHPo6Yn8x7VGENk6XWHPsPKh2FZU5UlOqaiK0aMHm54l0OP
4b7TtS1bNZdbEgv5d4b814kqfp5EE3r1YDWE73byIJ/sjqd/rCzjomoLxLxyfE8+
0jqIArKBD1qqx2R3/n9U5WdkRKQOXp+oLZ+rCKKz4yFIU5kfofnpI7yrueLztsXq
fULotvAmxr8Je3eYZJLp4f+sD7ddpJ21qtn5CC1CXWJ0GAY5N7D3rw1jtIi4LKyy
IcA/7Q1k2zJjjQLETGT1DZ4SPHPPEZRkVDzfmNDgJQmZ0jv9hF/UdW15YINDmdc9
i4no5rqwczWskkNBP4Kh+brw53V8NO9rS5OmoA2TdAS4PHcYxhTphHYOko+xqzJa
iFcCXo9NuiHyfSTcDxLh4SOA4CDq+OFx6hdgZA2nstnXBzS1z8hvWNUtChIHz1qR
vQHKcT+Ps12WtAwIj/ybjHCJepL+1ejPywtAOy0Fz8+qw+KIwledpp8aB9Abib6p
3W75OT5uPQqXlfeKVA4PBN1eModGmd5xOemdv2NLorXEpKvGMuJvxJ7wzzDOISNr
m3IN08Y55WJYzeMUiwxxeGEn7vy/9De8cP8wyjR6KAsnD0f7XAVFqtkXEmhZnOTM
Aupauifl2f7yMFL4SAY4uTOaSe1KvHKVlMDXl8XftDIZY8bu7oBaDsJ+95EO1XL4
Tqjs4xQMja/tmNgdwHg6MIsvObfXlEIuqJMXE6UvnxzAvFoVkcL0VdW1iBApjTDn
+BciHb3LAhXw1SWtMv8TjPtWB+J91qyX8GOabjig5p2o5GZIrsX7JrChXFOGm307
rbl4rx38Sb8LyFXqNb5ualBw7iN0fDhLud5M3v1PufFuR2D+PYs7mfXC9t6LNDZa
9uNdak0VrbjgcXy95gdPyc7eYhfiuVrRnjJhlPuhnQHOthBzEoAwvwPDE3qDlB0N
Kh5uo3uBlt3c54rPj9FeLxNwBBwJ7WduRbChXSM6e7m8ORKISDAyYesMXJc/P5t1
SwzK+FXuMkGxvuhewsWwjBNYlNdVVwPc1Ktx3AtS2Zj7j/tl89yyFFP1CM09xQoP
ONt64/AAg8jj8rq/uGnku13hRqTYjeErGIHQfMdOFEzbZR1sTTjjLZz3e3rN5m4H
LjeH3nFGAIj/meS+7kQ6IximXmyoGr4Gw7doSvIyi4IzpQ+WN3jIZEWhjDT4csyw
uMwwGmBGyAP27IKydt3E1JSWpEziLGYH2b+0/Yk/n42jRwn6loxqf7a8KnGWKQ94
Z/JM/VwC0VIbfXcNL/AISmvu33iW75I8Do+cByY7MZLmi0Rj33UntdKRbeVOsrm6
grMrO1E2DnWE22C3FmDiUvfw8EpScC49fB/C6Zs7RtS4WsX3PjEJ25cclUVuDjOf
nPmKN5pHdMVF5ENx8w+UFGTClHhupnQFbdc2e8dYTIIcLA89lL8KzYlJKOftcGIi
fvVSq6yXAm486loGsII1+PEKr8DasRqsNB4AKewfGjXV/O4zUG8WIBgBfLLWh3I1
j+sDyQ0HCR8aLrVsX0z0yerd8atyKCxuKFb3ipjjvrAo50LPYr59ZY3rRRiCu+pf
N63KCIbUb1Df/sIiCBZtGtutcfKFxHB7KcZ63yOvvVLDy+DYwXP8jeO6uzv6CrSj
5VHwPe4K/rbQEQt1qGnp+2+VMj1U41B4U1o1mTFk4a7zFbyrgujVnvPJchGzaQdr
AJwVarsFmC0+R/eju0zgLr0hdUkwFJtr8chn25ZF1sGih8jPuA3GM6nU6X+lGkiv
Uuc+htcG1Dw3RJ6RwoAUc/As45+nnevG0hNid3z98Nu+Y4+TFsFzQY2pk1PXME8v
m6C9xVJn1w7IFaQAjyNzZVZv99LvhlaonWKTttoA2CjQlF3X+JeM/KtsRatbX6OX
fK2Hu83fPg2akhtA0GasTY29Egmiq02B9jUWxJum7StU6A5tl88Opc/DauQJpqiM
nAVtayCyrD3ynpuHJLxGVv23thUUpbkaZMOr6ue4IkYf9DkBNVQJ3l+ZStlKsRmt
nnTP6fCur6JoE9s6Q7JMUs9Yel1p/MnkfFS8IXtohhpm3cTe/goEvC1gOmrM0Qp5
Pwj3Yg5gp/Uyu7cSE6jmP76PhRecK5VPclpZkMgwUxnx5dXXfuUI0837MWrT7rKo
hbRIgMiWgCuU4tyBM1AfRDuMnECVUT/dU0Qs+2+u4V40PmTzfeAmo+Nwz7EDiHXg
yZkIFnTYh7BD8KXJpy5WQNkQY2VQzmuD94qk+8Ll1P1DeqGBpZYWS1sLm3rxonum
pqJsyP82QkNpZN8mMj76LggxXSlYc8Ou2hkJ6vcglbdeTiLbY4rg3dhmEvn1ynWB
ny+piwYFsp7v9JdbnuUXc4kwAhuZMsdIV1bmuZCp8C+9PzRwCz/4wVl28tuRzZuW
uNZ+xbWaCvbYDO2MD2MqPNvtR4Plf9wBXWSHMvyw2XsnQxHp418dB9VfI2IDOLeX
Yqmp2KA1GD8THfXDMyZ302L5RDwhM9FZgF9ZN8nNE0iL0mSSO+uQFNTfhK17vzSE
GgLm3sMAlwtPJ6u34P+DZzdv7JfkPQvVPRc21OSsqYH7fVvIcBL87/YjC+/ltjok
QoqWh5u6coEDNfxeDJnjPWbbuc7zmyajzEgrGlmfGOr9wYvgRF0i8FgJ1MzTrzkz
zEX+4D1bbDp1F1V6RY68kS0XoplZYBLMDcFSiCzkxUy5x5JHLTLmKJnYCE485tSD
sP3CyDYtUqaxMV101264e4mFQpik2GWIfBQHS15MrUdtpSiq0M18iNwx9VMRYA8Y
s1pd/Bc81zo/hy8spGF2jUdK4PBezBVdjjMcvjRg4GGqTEqvNqSceB7/5kDzwgE+
oKglONQrn5SyoxPWTEgg378+uhjg4FvyoUmzZ3VW6Cw45hyhPpQUj0w6ENvGxaIw
m/7gZnktAIW3HVkhr20HoHUMXt4jKn5Wz+17pZvk7woSl5zGkFAftRW+iqwEvVwp
SyNflgEKGCDE9BMDaVC3hMG5E2tFeQ3XYFbCYKyELyiHCPb2XfoKAWGoGOcyYtfd
yhleXguQ5ouEnY1Uyun1v/0uUwcPzpqag8dcvsHBcKlgpCwFnu0T5HpLhGrajddj
/prir1mR4QWLFx9/a/CeOcgAjAJD6lKbVTGsUlUq2DAOB82PO0etVbdCrL47qxBk
fFr17UHEUabTb3gk658FZRsgKhUWxyCazx8mVxpRnX23lTJzslHw5WGIcgkf/orM
JaekKn1s1seyG6sEt7wIX0fU8f6vqG//X1u/Q7z6uHsENXkWToSSNvM7ojoorbMO
Hj7sWRIi7xN+WKe6N6ez4cLDJkzzuVfsDEwdzy+3XLL8DwCoCtNEAo0VLcaBTOla
eMOcXnNyslu8g+/X2XorrZfejnv6/atgzyv/K9R41OorYUfzbOXhUdcft5vs1wOP
MhIn2bpHNYpXqEAC/EP20HauVWhY7lRUIEkm7rQgBwiCq7PoauC+ITJRlglOChUR
TLlpP35/Rbsjn/Qv67DOOGv4WgHz525ZTcxXkhR63puDFunez2wGep/XzLkStTr1
X8fuSp0TZY/E4FgxdQ3eVIawUdPg6kFj4XWoxo/dkLc9NudTplE1mqJo0UazfWwo
rv9J1PFo4iMMP6JayMZOW258ayQ8weBVop+2yIlvyN2REvCHsTCAq8cYCdzn6Mjk
86negKFtlN3VReZYiq9fZc1ZuKo8vYKZLVM9/aLPGfW8Kz86MKUAkzecSnGHIIBn
al8gRKHc7tql0YnJaMAsWOIS2sXyeOJ5+m59k7tVbeBXWMb45RZZpVcxtE/nsXMv
owvPJebODDi9W+XHOdoJNornwbSQ5aj/qo6FxpdiW5xdWh0pMZ+2ybHDDzBSZ/iB
hwpgaNdajtm1b+9YKuxAo17nqJfVzuXFgP4h7s6Ud5ujQivfFlNjksn/rw6PFt+1
3OPVO878AjKCUMpQCLTIPiW1D+ywrjl84SRR53hLY3rAThRmPt5WXawjonw0R4Cx
ePc3TUzK2OuoYVvyZRzBdmmAM4YE2BVbQSarD8b5ofZRKB7XLiCTBYBXWUDswfhH
XgPRdSIhlEwfnDzT//Xr+lGHe/qNDE1QEIeMEenpOmLXSPHolZsXO+K1pDYnZi0v
2TT/3ushJDPqBvSsB7EQRMZ77O76mSrqDTtquvftFaH70jafrHAUhp18Cyw2UnAe
mM7iCAUMtS9yS4WEhF5puKl60QqQ+VC9JZ6WlP2j7Hsyy56fzefY7/H1aw7hV6Ub
u6+NPhqNLFPBiJ2LnWfKRIlnfd1IycWhTj8Wa0imACKF9A0N75XtR9tzb6lg7M5X
pLIWszhXp1SpQv5e7vzYOndRGJz661xtTbgAh1+czwW6EU2S0Vpch5oA7XdB5M9z
fgmmT909bvk4Jj/TB+pt0SSikTUtoZZFWXouBQdvijfU9VRu7hq6G6IGeBlSZeUb
+Hcr5KE+i1tHb9yfGxE6wJx3/DYSxfZo0CmVY+3mY5/19tYKEqEDYZtR7thb3hLf
VfiHffD+uccikTkkZi91TCB8Cyo0VrLvK+CuJ50saLGLl/dsyWWsRVVVG2hT7AV8
GrUOpbUSm77EYrMRIWcDcQBeMvLZqUVqhUsYKXlK8sQnHCBqdVbKQmegAPp1yxqY
dCOdooE0HwYhsesirMNqM/6BnRD9yPcyma5g1XQ9APKxdl/PNHryg0MztSa4qWaB
5KVdFHiHfn0FRqZtGZNW0d+EIkczOIYQmt0ot34xru0dDZGPFaIu7qmIAsC2pNmO
nDqbf6UGmh5rA0+G8DKatyONNLLnL1N2XJTdaoiygAki7B6bXZst0gjoMtX0PnW3
O3BJbCnfGtTSKfiWewe6PseYDC/zmKgKCYZzvnJ8aB8trkF/He+yX6OtcVP4SxWz
c2L3RwRJw//ca4KhNDeWcWcS2RI4OWM8UFGatbo61AOqRiqFhggJp6kQOOPyf2kt
eTF3Ktka7vVwXq37COwDznXFRMJn0F9WYzX3AjVhYtgwVA6Q393v2L+eSVdloqhQ
l6uu21cAHyVpUOJNYf6Za8MqotIbEkZYmZ1WGByBQCDyObgINyuMM8BgMvnmzSqA
2TbDf4QHkx18Gl5N70HQh1zhDhPploL23nx2l7Dbb3hnIatgM3ZMyfgZ0eCpn6Tg
PYI7mjFC7iINczuGN3zImgepDTAp0oLW00PxI4CJjsd0R6ZzqC9iribzUHhcfRls
2atvSTNqEARozTvMGilIvO6tBjo9HpKvgmAF/LCii48vXAsWDfXxtuALcg4SuscP
dCDSWDJb1p2UH+E8CnSVlBhE2q12N/OGjFOJHYTw/kEXV45ay4pqWcHvBsNiA3z0
+Qm4NlVWSsOsfKbL6CFhU6S7Lqy6lKRT0aJqQW6yYg/dwsrHM71uLOCxj+i6kGk2
UTDlDFRlh299VQ+VXhzA1MpnOb00vuuQ00m3WAiBb+xEy6NJow0TlV2WURwnkoKw
bT5Yf6rC1jE2kNJhwGe50xvYZDXwV82t9yLz4d6tRFpj1oMRjfwVBpw2rb3HRMT3
HRVZcWcs2pcxQqRPTiqOfrfCnkMenTg0CIFiqxoeluoynEUko85Iq3q0J/J9yTv1
L0VcPYLnQVMuas+Eal2wqXcRVYYyZFBXW/CFktZtHvgphbY94rlPcY6NJIEv/0UV
cdboBKxI/smX4Gx3jnpSXVwShX7RncwB0LZg6kqHJ848okDXV9qqiXav8dhm3kEY
MxmW/ngKpcHArUEJFNpNPu1gjjbYNncmWTU38sURDa8dJFLWcCLq6CxGzKMjw7Ez
tIwuOvT4KUi1+wCYSyfRU5zFsMSNfl4UmeufGMVE34niyoj7kenv7OU89nPGdQ5L
jKoeHeWNVja4722MZzLLx94ymqekBtUR1e6jLK0+lYCkPHcIwacntpXjtVnttIgR
r2k774T6d1/QdpQSzogP30UQUDX3sB3uHNjFmvEvbuBqIAmz/jSB3AjTahSncGIW
zINvKvn+d4f4T6j74aLpc0VGoUd3HroEIaJ7uXZberfNZKqHqF9MIpIZqpTgr4DW
d0ENoHz365AZYnRYoCGydqbiL8FZ4pTEgVuuNWXT8OXF6sEHz3cs6PJuKoYhUgsq
V0vjiMCaoUFq3w35jDR7EPc1+9HeOQ0RDxOlZ5jbR6zMyaV+CCrrgmLcajN/z9d1
F0P7xoMomrlGnw8+FitziypBEq5RGIgJuNlquut9khLbJZhxnyiYNx/9KOZL90Lx
wQScn8WRPtoZwQK/7K5fU+QjVrFelVEm4P07avo9iWRWCq2RP2zqkqr4Ox2/c/d/
m6lt2pII42DyxMQ10y4bX0KNvRNcmsH/qlGTgX38dAh3KOLBrMxIhWmMtp92IoPD
M4BPGs/8qg+iBjLgSbZx5iyMSWLTqBQPM9NgfvPkE7jdNOSwE1CZgIc55S6UlkDu
AIq7719HYpm4e3Bvo7nIeREh7yeQEZco/rYEZ9Akc6/uXAqpMFrws2NUhlxsMnhs
ZjN4OZ7jCi/gu837zTE0TjXc9hg4MhIhihWZ/Px3hHI736TWuWN3INCLyvMPnmko
56s5pbHuevsabHb2T0A7Hxx2b4S19uS+NG4XrD97RxMVOwAbmk5u2sadR+Vr02n/
tu+jkjPy2+uPFqGNDqdnneIZrysgtQfov/LX4RoTAoXv1R0a6BclM9liEJIHKOEV
S/ZGg8mczW3ADBXzlBQmP1VGbNd/mTldqQD/DF5hjqQkrXWc0nrTtX4822AthMK6
/LFmbepTkXFOpndXtIBzEQHyrQ8mD8A1zjeMquokuKlSz8rucCJ1ATVVVP5KqinH
QIx/YM3b0RMwdnDRRt2M3Fq62O22lnj7ZFjUiPnSOojUoWRZa/BaZnhblhW5UXLh
gkbu8YCYjXqcAgemcocFo5zyk0o/PnD2A6KviPo0PAfNXbrB7Pc5cyJLWaTPIxqv
SuqrFJtbK1MzLyFipsX4q6OgwLD0dLwIDQVp5Rdy5SPABPkR3tLutq95EXquSLvq
MM4+ASYTvlYGVEVkzXS38euXe3X7rHODhbIaieov2XG2UUqIhAfYNv4vu4xNV/cZ
3j/oBEC0decyzZKqpRM74FjS3HiJTqScrVCJCVYmgSLCnSfMvVH/x8cebZtxiFIo
qVseBfBeRDPoZO9VkuGf5n9XJeft5+xBGgKQWiWqCo8H3Cy0McBLzXDDx4zqRnsr
3bO5tJLBKze9fQ3pngnsG3uAKaZGPLP4zNFuAO3NZB2aMUDNYi6HjMXKirhjcYi5
w+beLa1/VmOvXt9FNADeAbYRkhAO1ZUnqcGmZUQ7vr9idI5y9a6yaQ0gPFtIxNN6
ymuJf5MEckEkwc/ERyVRkEzobXOYzAwyTMy0OTCRwbgObPLi7JWlQrGPiDRL2rPc
5hmDR1O/T6gCRt8zmOqECIiSEjQVfFhQPfCqaoMHfluspr00xY7OHuGdOLKZwI9a
qUj9wWWnJYSf6OxT1Ns3YAvL9gSq4g51zMPElzx3fAbI0bf6khxmCStdN89gEGFU
UIt7M03TDtkEq6c27BNV4y2NrHOpqbDiQv1xMmIiAoJGSGkXdCyj2TeeKW4Z8WIR
mwW6pDyXpCggCoKb2u4PY3KZi4JDAOiLgHnCwHERIx0H+TP4222DcZbZIm635hjZ
N6upKRDHmkl6jSL8DgNEW/e5A9N2sphHGRLTHmJxdNu5XROHXPHzHlK2BCvPLQe0
IX3UK2FZL/HbOgf/nqC0EWvGKqOdxU8GzunzDNYZooMkhoEz0EbrjdA1Cvo4deto
151rqVvQvVRcw5XjusGgfHvt6OdpHEQ7k0SWeRKMjGZgY3uCy9ehtJDXWUdFdE+k
GyLi+E52X9Tq+IoPlJmdKE+pGSQmWEinUspMyZOlJGJ2OhclyUDdnmfujGWEqBOH
LiS+jB/qM5m3cxavmfniUkg9wcSsyRQlP7V0jQBKWeq1LdtuUITFzq+/U5a5Hov3
em8FamUDKoscgVJClIVsQCNqnIP/KtBKfVD845+U24+Nw3BQuuQdiQPTNX+Thr1H
xOLOizJmBu9s93s1aaaKL1nj7cLyXkfSgzCrgo3VPm7MW6RWRiOYRIwMgUCL9ja/
654LysPCqSHtq5Cp8ZuwOVaQStyTRWFfXzwYgDo5+A+7PVVUDgu8qxOLarORkgdt
aY++ega8q8m3q792v6lIAM6vZj/LDro2qsW1Cwn75w5bq4+NA1RM+01eVlmYGIrh
6bEObIfS1BRUOaLPfHI6ka67cleRPUcUGXwSd5yHZ8P+uk3Z21esxWd1uy5b4gK6
m9unpbjDN/W+6yUT3BB+l2oM6eGGdUS9YpVkSM9y6CI2B2l9t7HKxD+5KKRVjbld
wWKvGD4/3YeGvlA3Ps2pEYFXngG2mfPIPI6BUtHvN9+/ebGJSZE/b5Vvvfr9c0Qa
/fDCsGOcr6DNktV/DdtaNOlfYw1OWq3oTr5OYmsgFdlbOE/Sc8RgOHMa1y2JU6eb
AnHHrN5zx23cu0SrmATfXg/5KfZ599J67iiEz7Q09Ne3hG32zcoqcjFU2+/abIVR
89DW+YaDs041R2SCkLATbh6YjEVUazajb1utsjw17zeFPgJGaTN3l94bG2bNSCqm
q9ZwRzn3R/Za8GVUpA3tlGkwE/JJTtOwXsVhA+x5fE7pL7cm4ZNyPOXUIXOqwHeb
NV6FbicHjxn4WULjF0ZCOnx8twkVHN05w9MmWkh9t0lzfGn7njPu2rivUNvO2Bgo
gERmlSerxB/NLqsVTIA62iK2/rzDPRDXRVocTNpONQZkr27UvpN+7JaV2u4Mchke
FJGdoR52bn+Eoup8fE8dJfV3EnkcbCAt/Emsb4rqnbK3sMqpyiQfjIh5OgmFc3PF
GLHQ+oL3nKJuwOzAEszoVbWGUyKMVINOGxeTnF+iLlmIQl4iJ+G3S2pEsbOsOvJL
Rho9jsfBU/1PMUP72UeEycQVX8IVU0CfHlqrBEaaBv4rgoTGK550Vld7XAixi4ra
iJuviubF8Aytbx1X86PDg+s3pZKxqVfgkAbT107xbZoqApQI/msA9GnMeBYKyCFj
yIXeimB9yRw81z6S+zSkN1huC1ZUea+uQ6nQqU7X92OcKvW887uAR3QiYl9g7IAd
cwAnoQtCZrURB96PcgLlZ2mt6YwCrJVeWFdEIpJr/HJm4akZj1mejS80bvAVhJRJ
xuIpftNULzMzJZns38IK7IZlGdfXYPLeD6Up0xPrTlLejzbWQGm2/2YkjryiSY47
tr7EddJxJorAzLtxb6BdB4g7UdvGNG9cxBiG4dJri/hiyPP86fjSjUfNxfTFnO9O
7KKqZPEwsPzsIacaPHfTqD9p9NotjgRg31hN2BRs1uX4rzAltcVWBLueMQUpWPie
jCJWVrSL6RWeKi97BPvjrD/rTrQthl5cHfcE587JuP5Z697+oCAdIK0lF95x/dWe
JksnZ/mzGWUs0n3MN8k9CCnVTFh+YtWQMW5vFlFTc6yzRXwuRU/jB+ANPaOm/RQW
GHSs4oFSWv7cXRrZMS7ru8+pJgzl41XoS37678de/k1YbIJNKK1pIe5A4Z3bcn7p
a0zxqjJiyWPl7PdMjvQ51+J7TbdXz6KDEh8uuqfCqb1B+mp90STk7CzIojESljYr
/o51qB7LwnusJm2CLpO5EEPp0b2Aw9oyYT5UDx2nhq5/mToUZUz5tp6aQCQxu8+O
A3hrMYeO4gP3IfBRbwHApwi8ucAmC2u/0WnNusHWn5StbwAuXdS1SKWb3AjlochM
Hf6PnpAlw6OejVvgX25+QCkdjcBaTTzfyYqgCFzMDAq3emVscBrqXd1Yw8aZbO+k
j/e65MqJs6PKCItDzfFiblUeGGDE7U5WbYOBxsjuQrF1nFi36Zk6hIDI/4ACRMmd
QFc2++RnxP0hYH2L/a6j8ZAXXDcwDfkzEowASmyhd4WkjQ8tbiVWut9rdycGdtLk
gt8TgPkDXC6BZlqCj0OLKAXx6d8M1FvMyPQLt1RmmIF8ITonV5rbTfup2L8p/ZJW
b+vZzY8mKKrD0DvaGhcyt0Bg/Cm2zLHxrUFZuUE8Dnrl4DyKZJEjNJT13VM55gaM
+4/AfiasSKo5TupgvV3Vrp5Eh4RNrxwVcqA/4BoBHmX1oMluItF70fpLBs8h2cDQ
WPr+LnCggJ7CSNk0lNFWtvZdWx5Z/hQqwuAnhNGnuoGgQ8RUXxalrxAM0tB4plJh
fTiyj9No5Mwv+nQVAHrUSuVkmJhOWtzGIEDN1anR5S2tcwnKC+aJAL8lus1VFDNp
oB2x+UaVFQRI9Whn4R/tNNrnDKBYqQChhFUkmvNc6hccIk68/iU0ycrotVSYuToR
lGVNN9qhbQFQI1YQU+zLroVBDkpfRYSWxHsEVY7j17RdjXHj1OMYPWJcAnRcVA9O
J0Zh6OpUch/Y+baNGbGxw9XAquv436MHEQBxuS+HD9a6agjZSJtLJ+V4oBJ6lvhV
frN1/JhC3KjciFJrzScG7GnbPV9AJIQ7ttTH3zimMMut4cACLto4EwHQiTg3iygf
7+nJ8mUGhPE028NCfLhTaZupfeOYFoRi7DMRRJBiR15GWrrobGdDDDm5xBNeM5Q4
QRjaa37ipgz4Sy7BDlsmDo19N8skfuI37Eir8cUS5jjp/rAYFLEUnT7xIQtjAXbe
87KcvQ5N3ee4nqY51b6KcOhB1zbh62IIMc7knRBRI7hG3LOF+5crGww1zEJd3GfX
Vp8NgMbXZ/FCT2YJYnH7/jbd5c4hgnvWGWVjScIvWrSgywjDWbXgcJm7zMUn2RYx
rWrxPM8RtznD4FmLNLyGMQmNrd4j8SwYVozlYWBSlkHfE6KCfc+gtQ+cKA/PIqVf
OGSJaGE5Tg9s7qroDNzSQnveVX7EACBeKhDtt+DbfGPsvxJsV1AugHVuQPRhjXVm
Ears1l5vat/upprYVK20DjCfa1m5noBEVXg2qMpP7wRfH1WPTARfUgXe26lhOla+
ir1Iv2WRjx0OBUIJqwrJC+AMLR15fiIKtCqRu7XVHVbCw98yohjzEdoAthK9uwjS
ZPQpihAvpi+WcIwhv33yYjzqpUUcVPfqPdigorN2AxT0UFJqyAzRgWtXV7E/VKsy
FPd3vQ1a9fxoHz/htKrlFTglRy65OIdFs7f6Lyms1hYfTvF5LBWs4agyEZu6liVk
x77hY92Q6UjzZQ0moUTsSuc/PXG1TqI1ccrss2ZqjBoXyGoBHOG9/E8ruA9poGei
nWiKOJN5bVUNQqrE4WCYTgwPjoncqtTllpYH2DpWzpxxC8IlFC3JHiR6dFUBBWvw
y868t7ukQjXVIaUhsCqH+I4auRUhTkqwPFmXPfGIr0HL6k9MxZlzJwvpg4iLs49E
BbpUqHV+BPUIyy5+vho/ZJk3PGJ5xP9rYZGOmxyiDxZmgvmZj1ZXCTChRaOZmpq6
F7cyogRmC4xnhsgHK6F1bMjG0MLOsbOz1YBmqL15BzHeb4Trl5nG3EPrPhYygpnd
NRWhALsXd94+P0NTn4U1z5OR1Nysjp45tNgYqFGBRzVOCiv/wH8V5M20f9edt/WE
VpoAtAU50n+uIEmPVbGWRgxPxViXK8DCDDTJI7Rsw1Caw/7OkhE1HL6MSq1+5bGM
TIK1YPSq5xmFPQhjqr5LMZlSNIYIvMNmtZFyPCdsAS08IHS+4nsCOxw2mk2tzWw0
UosykYFM6Zvk/pRRPrhChph9edRGyRgyNr9gHrw0hwbJ8Zxh+p/OX321QiovINkd
fLBTCkwdUd4nYIBRfaRbPdFGD8u0+ZWqivx5l4d8urZEKw64knlBWD8Vf1xzr2Es
5ENDwuZRBjl6GtnExWIP3fPRRh1fBq+3LiaaWi5S8J5bb2SLG6Lq0zblftz2+rr2
YyQ749sRu6HgioN7etqCWVb1nwJpMq9TOS3rA+DoypPi2OWsEm9TZltP2RQK+scs
PkDqwkNWPOQj/d3D8kw8Xo8NSSrX24zg5tdGGbXJOiVGmmHVO8qcoPhggHCEjXgL
Kk5i2UN9OZcW5SqJxiJeMpVsJZZy4JzMFNchetPjRc/RQM0wCn7Ug7PfWcgqNwKN
tGX1x4Zvrjph8pYSTXdebETQFxSpDxZddvo0YzIfrgDKI4yTGv0MDEmHxzzQJSRK
soJ8RKksYomKgZjoJo8l06Lv3+yB0ZxZArqQCZ/ZBMPNd26HxM7OjXYdE5j/qc5O
JHfA+bEPiG0fK6wT8LXr1jYQousikdcnQOhiPrmKrjIKUzW2RpiKd5pNxhmqorm9
OJbpk1l33EMQgxu35GLgix51PKaAIgSnAPNDbYjHqPficwFOzzqRY8Zuj1ehFGCQ
mebwtGRRk65S54wOwV3p/v4F45HLTFVMiIj4NBJ50PZ0DJGpzBNY2m2IhuJt1OIL
aXzEQaNG+H33D8kGd35szflZhI7IKbtdev6uvQr6sWlTwL7sXIApPyBsawhXLYJi
bzrvlMEs18YQW3mpB/n9CkGg/hguScz7XTNOU8kvlJf7LbOdlrz0KwV3BkavVUF4
9k5ggVDM5HMSnC9km5CATVQ04QmQBjl/IUgaf09wE6QKPZwPMPbKKOPWcwbhl8UR
3692QaeWfTBVOTWsOCClv6xI1h+NE9Qc3NWLnbbvHdeQ1u88kLEF5ChqqrGSlzjn
sTNjM4EJ+iMskjMA5OsZwF/Oct0zArLTy82JnvfCQ2jCG2J0V0mfeGatVo/lYBlU
SH8yArCs0hgizkidFyQfM9FykYW3znOE4R8CqbXoMdZYjjqy1J1/A9nXDF/gfR1r
7U1zv1HYi7Ac/CgZVMDqYFOEQn/kUk6U6/+WH6XnSgpcYXN4aHK93X3iDeg7007O
ia6bzUQfHpIbOuUEhQn09mdDSUaj+MhhccRKVqsZ40ZfMdojGwoqY+0Y4KGvrhzn
ZDr9FbjEIbNwx9bUcLW88ZbzkrVoaOSQc+se4lL5y5HEY6Jo3SlixhrqXsfmwtfd
wX79qr+3dfyNSadqCOjeiX5Td9omjn5My/q7qp8O6M42ysm8BG0LsnCAkBT1/XvJ
zBaISoBARLrAvZWbhejORSJA7uTYt2sauUTVUrglf24jNk/yW1WKz5AtuIqQOXRF
iQ6Ckfjxtn2v79S5mmdiIqSKZsaFDZ05aVBY1lQoN3jFOJc41jIHKz9JQYiKtyhp
wGul+txhasanSCLGaFxCJNLEjek8NOMq8zoPYbruPe4DtHRPsR69X5h+BdGbSPbv
ydIkEUeCG8jISivCfEjuYxD7coP3lZvKmndjFQquHClIKfYggACKc19yZ8aI839Y
ZXFAyroOHtRXZFdnrXI2Vh0KZvQpEEG3vZSRApWu+9u83QMwLb48mYwHa7MjUCrv
SvzCaJ8XdT1is1yUw5+JLBarwmhfgOI7vTJvtzQI6lIRrZDTAbQxjMHE/jY2iJuK
XW9CwNw0aaqjQj9ssfNxiqYUKY1rVUcXVN+wUvfKB+LCKlIMn0GGOdG4xLYCEz3g
CrN4Jqou2N79hvZzlQHU+ZPxXLREVPZjh4dDcFCfFhYvDsKH3XjcT1fX2Ql0mpey
b/9sIfFdVuN7eUlUgwKHHzoP0ZPUPvSL/bmx6xHo/TUyiykrGB3S7e/ZVCHeJcsL
Mvi23Ge+9BKZve3F8vcy5eFIjyOe0ETgs/aKqe7qF4hyLDLJjbCS2fDOHYHoVzJK
6uJomWAY82Wzgo+FXoZS9fqZ759iv8vNsW1jUpBC6F+4lgzXobXHxfkSgzavPhn6
VqPopDKQUeB2qg2+JSa5U3L/kO5UD/DjcV/eBl/bMwWNl+WA/Fu3ryDBg0N9Hmlt
+BLCprZEB8k+DN3hOnSkb9CRtUWv3eQ5XdTqR+gXCUiPiHP6TWFUYyOafjXvhljy
gOCM2WHikcxm4If8bJE6nRsUEjqFjk5iO/EnpV1mvPClltO2+zKhGjOHsNwW/vqy
zc+T3BXHUn/KD8au2S99V7t9W8cHZyAqiyRMCfef5ZkNEoLhyZmwAZlAeof7qtf3
KBPoYddNblA+HYfU/TGascSI5WV8oUM3PxayW08dmUxZTrTctgHiM3LRW0HD6R16
gvgT97CSGUMQOBCsVBXSHzDzu5AyCaxoANxSRye+cy+Wuy0wBeFBnYjaX9K3iET7
ig58pEeoHmak7IiygoHP+Sk6ul2l+wIfB+aunzALFg+ZMy+sOLPvmu572zJGkSGL
UfZUaSfSMj32s34r0vIoo3XjjBmzN5SDO/sguTMHpHcIDNVj2PgzQItu4OFpnKEZ
sUl1+MBtQgtp+DQpwmPnLSd5Ygd9ByxNBPzBvIm0R1t6/FK7NTbvYbvuOZX6nkuO
B3grxgQtA/o+40i5ZWm/jFOCqXYKYqXQ4VvW70VSlqPzFc02zrTBxOC5YraLzZXq
LNJApDwD4483onQtF+TKL5EUn7o8DWZwsCVJUO5Gn715zOwtXSGDKL89l4VxRmIa
B8VvMGcbIKeMS/v/uRlyRWCZohHrvUqUOJuqDvFREJIAHydXxiRHcdDJlcO8iwYV
wmwj3BIKApnHr1zJqEnyePXOCGMtkx5GGe+E71PN1O4KVQxqEO3U66PXWdAxge1O
GuT1SvQNOvwLz3p6v4MD97ussjOfy1aqafLsZrcDI4Y4PVDOAwIzJS/PPmObG+aP
rhcaNLMwZYyEyM9pBwmX8f1WT0h3cNSOR/LHBch/tRjoCMwZIinSxWeRTJlYWdl0
rpPqM4M2cWKlnL3hFM4ZQOCjDeZBxcHrLCm7A7yN9qFIV5xcQ05LAQXE4ufkol+X
EpbrEtR7z6StUsNCnjQyfYs9hVERHuHlz+GH84LxL3dHVT5r3pyjI2mQM32Euck3
sB4Kk/bJT5UDNKbnp8/CsuIxKXOvqDGrbfL8BZtsh1ugJnkTJ4iJ6fbynS9RrqLO
sc1wI7tFiaODYBwqO95kKv1v3ZY5cCGzTIb1NTbhoQrIba1LIodtPoX4wNhd84uQ
jXSPSfexPVshKJJ6HckHh2volYG+jGyg2hVSEcUwjBcr++bjJe/faaaaV8nsO3ZT
cnpqFPpEABGueobDfc8jfNSjsewJSge7zl/jHybGsMklw3f3Vzf6gXHHIJIXHWIg
BznwN62tPzqhD5nAhCYLzdae7uJLUz03k/uIdBnVlkcxJRWXtUqUDrXAz/LgvPrf
+pI10PTGE4OUsWCl0o5aR+L9wMC8JBCWnVrdsWOFH01AzD5204OQQmZmqmWfGhzb
ZfVXGV6LLZaaLlt0Xz1rkNA5FEbrcyx6M4TGOqjC70zKKukn3NHKF1xJh/BJa96E
POiaewnnT97M7rgXVICQfj5P28ARqXsYK8ttfKAszs1JbpeIuq8fm/2Z/gh5c0Id
ZKDs+nGK+HX9x2MFFdznD2//9uYRvqHQuKalPUsbllYg4ae9cOGyc3/uk2Qzy1d2
ZQ8ptDJ95SeSUHu8+lY/NgfowtBYj/Y4MzuDAvBDB3l4LYuNqqTsj1W9t1jut+XS
OLkLCeWoloVw1sVlUGJGRhBBbVPCPcd112d8ECfF53kVpAO2C4tJLIrnLricxPXw
4PyMEVCJpxzqsxTV32DGIR8FDPeET9I2wUrUenYosBPNVQMkC2j74gnBc7lF75p8
Hn+4jYyZxK3zaC9ieJxnaAv67X6RgGH3eRWrgHl2L5CDb+brLs1P5SNwDWCcjs8B
TeC12fMVcNijjiy8XYVsLRm3SJW23xsH8SXHFL9nBz8afB/L4fnkQjRvaC4HRHSL
Nw8Vm2cejUknK70vEp1MPWcbpQTL1+6OpUSZCuQ96QEdU15V3ITM07b7zw23pA6Q
VXG4WFzbe0BCsYWTi3K5IcJqXjSbQF8tt54oi4+fEvT8i1WsKPZebYl54fN3zCwF
ABYFbyY20W7kumIoMdrF7BXabrcnBEIQZNuvgsn4U8Ndt4WoXItzwsVwq99C1DEB
SlhHlFyb+3v0b+Izu44KvdrTgk0NDuGm1eapJq9onZ2fKO7L0IIKN2VPXutb/b3I
mtFG7nX55oc6o8mFMfN0Diq252D9lkvCCC5tVg4BtkXyUEvOjpySZ8KNPG1/AMG7
EXhGpGZoyjyQYA+KrLfg1lANWiB/kFCn9/YA51vzXOSRhQbGOOEhfF3bIU6rUsLg
SKqMgaR+QtdFzC5+0a1ZD79e8NWun9IBFxa6RKFBFaHovlXO7F2ipA7dBE2TkNkN
ZqvX1b5XDnZJkO2n8ZAyEXUEtso2iPPQetru9fCuSiTvs+1KsYrIkt7GTvzWFb66
DRz3mA/JFupffMYXGnYbFsU5t9Fb+I/xbyBc1rwa+gs9YGjmIC0kLloo3rzScGBp
AXREWTab/699VDrMtBLPXuQR+kXLArwyZGECQvrIwZGyZXh8QNxARIB9Z+Lk+IQJ
XSF5QssGXwve+c04ZloCcsrDF2qGWALy1WPGIQQV8T0iUjjZWMwVu14w5qCN7bv+
9EFEOTJ4Sd2NbSqM+RoNnbfm3eSrDP7x77iw2zsLhHIgaHzyEOJUPFlRSUXegRhV
k6yL2d2qUK6P9YdJBeXNN9xLH3YpprorDNk0SN/Ub3tGVM3rZGpEXFy5kS9XdA3n
QepXFVqbmbycsUEaQDwOvn2E2TBv9OSSWWVVVOJsUnAh5jwUKdn6RcK3UiZHRAaK
hPUemvSD5NE8p79G5p2Ztq8ct2DPCs0sQzl0AF2crpjks2BM2hEkMuIJrXSWWae5
vA28fmeDBN0wmC1vBsxF68dtPBx+wK3zbF2aakaiWplLORuDpGbb3i0SDGvmgdGQ
RWe61Jnym4BuJNjxmQNrrPLWiB3VeXvP+HeUbwjxgLPj61R9TIH3D10j55dEVZa0
i32xIbMxpjkiOYDfV3HCSTck9GIJAflmWu4NvAOTW6dHEziAQJaliWw0n3h5cIwH
PXSEEkf7/P2mnf/14ZKOjVcS828VmizKIGbxpKxKk373POAqNn6TsGrNHassjPJ/
UR/d9EGNMpLYqk4wHjo0fUXVmhwql+i3DGzPHL/CaBb2+rT47fTr4nzPis64TCN7
ulem99u6ViMcEycL/mX1LC5bbd12LWcrv7DaVCMmFh0QYOIW0OmnmBXGeZ2nSZjE
j+O4dazkJvdia/oecNFXqP+loC56vTihwxmzxkXfDtqNaQzRfhybmxR2jssgyQE6
y88dMk+xwkFnzNqoy0QWnmYvjQi3houxdhpSoP/zeYGfkE6DBQdmtyMbHfMWuFAF
Em0xn/5Uj8/mbXsX8E2KETWjvsKmV28Mas2gy/XvGGZ+rngjgCkF+UfXrLBdzBDS
vFOcQEC7b9u2KUUG9eAoP+4n38aiHR+D5D5CAKz05X8U9PQ/khnNlCdghBsdf0Ig
oGsnRhn/C4hsYh8jgcv/T8YNlqrYJpZVSLf5h8SuDcF8JoWok6dszwnRV1FxPUjD
vQhtVABd4twKOp63KqX0/+AadUc1Mor1VfzFs4gu0Y5JKimNcdZ1qmXMJ0M210pr
ajgc8ULqtQ2i9ejUGab8BCzyF6pBJZ/0+QMlrpc05XlHnn/T2aZpx0OiaVX+gsaF
H0vzs+4oe/ObstR3KnfxWGkL/J1/qPMulNRSyMw7TwGan0IdV5vK7PSlU7dbcm56
7eqAubV31pEUaN14LfP7v5uOudg3DzHyGXkQHYrgdbE9TERens0jIOp8S8YITIZw
E4p8EQNEI80qs56OZOX1h4uyuCPTTvu3s1CnLJYjpybO76fSu6/Kyt+Mdvjz1pOz
47W4P6FHnvwbT37f4lYzbf6LoFoBVkxP436N/2+ZuAmYQSQHwepEBwPxwAcUoqJH
4DvLE8HnQFoSRH7Z/YyKjbkogqQ2q/Nn+AjevGkf5ylP95din4U77A4kPaZ32p6e
d3mE6OZuwdS07BHd3aE6Igde5eNepPr05Y7ouDcvYZgKewzPtlornj8TD4ijsXbg
9mau9RtsvvTMuxNuMqjN+oNR13IuJD6SCEBGSdzyG/N6u5LS9G0PG3pgwNJMEkOX
IxKP9KF6BBwruE7pe2nTi39nnv0A63nMnigdYAOEDC9hsEkW+GwW/9GMnbWwIpCe
YhUOMAYuiqRVMTAYsZHKlovYRN9nulGNQl9TGvVdLKgRcrYUVKmCakHHF26YTYny
RfzbD4pOsMhj8FmZ5hL31iBGWtzGhaBnzgkggEMQ+vbMa0BwbQlhfSoQF3cMjRbq
THBGCxLU2t6Wve/SSYSykNI5UMLZ1vJWhyBYTA4Kav4p3Cv+Wgm9pUuPabfoyb/E
m3cU5rr3L5LhMU8BldTz/jeG8LXIjGRP/SfuHYDYD76yhUQQvFo43+ChYKZd7AoU
GZbrQDPDie7VdqgDL1MITzep7CMqoYfxs4VKo0p72+sr9VeGG05ytUSb2lJ5/QVf
ufyBOg6FBRMjEdLNBm6vAznKv9AAa7O/DWZiz0NaTNvNA/CcMQ7gZLhGz/FzopyB
QFzkWTFwarcMJqnSnBG6UYAVPw5FFKjV8a2WsywZNkb0cwnL7WvjDVStC7ld6M29
57zMQKs3E+MHfideUF0j8R0Iwh2T+lq9SzayFj8lvIOQLdoSS6vfW+enD2wmy5sB
/Z/rSCYXZ7XdXX9ehalVtxw/G0IoqGFTs+DGE7xQLhK2JMwIUskO91aKzA0XPjIj
b37S1FJMHV6cQsrBtf72p/BJySmIEXFMPGgKcr2xpICD5xXvXqOKgL93wPN/0klY
jxbrN97u7XJW9t6tg9vnG2BTu1xmTFUOKgFI79VaxLLX9Bj5l9nEt5DSEDNfztWl
F0uADxowTT98yeJuvleTkc9YOvjAVs5CI7LNDj1WJXMnqD90iiBbRsjCzcfoCQ+M
hBfELiW69IHj4slLoPolmlhJOxwRy3Ic7A4hoSJ+QP2O7tr+OX9Qy6Zuke8LvdCA
FENp6N02RjRWd4r5B+WgQHE/sZ8hP+0XqcALAcRdoL7gkkh/qype8omYnGlfln9V
iQ5Rm4VaL/pgS9fdZhWTDxapLbkGLVbkUZihCM5ECPrHtUaTZzVwS4IODBiyK5ad
4Dv9Vkkh1Agn5pAhd163FMM1TzFymXZ1NM3p3HZAMvvu8ASCShEbjHE0cAekUFFq
dvNZBvGZDHKfzQE7muKgWFbpIZsl7lLaOnaYEtdLnQQyCRBXrkrG7qskPmLzMbnA
nnJlvFySszamtUkp2E6NUOid6FOGTt/wutShrUp5n+rW+1LtFUEBOAsB3HlAFr5p
x04sG5oWFSCJ0OdKEgxlF+BG3Jexf5Lp8WEbHsSamC9ILzN3kpwHTBMdFBVUnhJd
eD1JD2tSyHwEYEqKQ0ImXbZ0q2s+GUlIzTxJQpmVYWmIHncY9FZHmfKWPjNOQZfE
K5iK5clBm6HFe+8k3NTsiCigJ/t7MVRO0cSVQkzGbw5Q9M+fS7qpxV5vV9rMTok+
Kf1Qqe9mNhEgx4ACLIvboC/KYrYSj7TvcRQtdQZmozOgpIkjnIATfAyFVXUuv8bz
L6bXTQ9o930fq79BZp79Dw8eaaiyAPIv7/j5bv6jXOQBDMMhR3IFsXqASsFbTPf3
BEfcUj2FXE2ataOnV9S039zW1imyQthzmoQGfXexne/GhfbGPlpQCIBt3ghYrAJy
nSfJoKtECQJ477+nMCBQ6c7hY5jhPSOYMrytEeZtfuyCfDU27HxyXphow0RkKOu2
4w5Jh744JvtxnWTqkzn9nWhkBSmG1ihZK6K3Fcz02Uq0KgjUEaHr38SUIWJkjzei
ARp/Q9yNk9A0MsLYybhxRNJRP3mPUA8VzkXjXI9r08BEC2hfPznXR4VfEYNCoy69
Ov5OjbG4+MqflO180Umsbp1ALjweVSZh9pXdDJkdmDzskFLMbXqbd9Y24QuJk40v
n63uEGPeGZsGXcd65LRVLQP5SCP569G0xiCF96S/mmkffvC6jLcnU8rSOadg20/3
E3ccmo89X7KwsYvrLR7fQuX3LHPsLkZbVBgGwS5rWWKrtiueEmtqeRYDOcWYwsyo
Rya/yF5XQQELJbrlwiAShvmt6I234Mmcgp9flrgNH+yfvUOcXn2Q/V9dIzUiH1Ob
vmDmQ6q4i49VwvyS7iZs2tWcRimWgSOFtItI8+2RudFkJHIzMFFpRSemEVDfAl4Y
cFHHY2dVZfIojHbdinvQO3VV1FWJcKXX5IpckGE7QI3g2F6W8QCZF76Jwtvz+iRN
dffmfHJgATctF1hufrzh6nUP67BqiUKhhE239PsKv+xvpQ/UvH8FioWS6TYi+PvV
R/9z3zgV9qpx3jYXzH0/Ffn0nGy2gF0l6E9V35hPn6q0phiQ7d82E9Om90khAYW/
PILw8/Z4zgXJ821sG9hZXKOFn/nIyR1HvMW0OI21iqBmANaJkjOhdhqot6H2Stc5
ew1NO0iS/oo0jn/0wW4HXMeP320TKR0GsoKyo/UtBL3xAIKxJGuSdYCT0bO6dE/w
vMXuPc8K9WKombkQVt581W2mKtNOZcerUnUecZ57PFNoHjrFCo3edM+p9yfvuTXf
Ul1OeNz2Sem+jxZfQ4MgTLqdfk329nkG0vsQexisN4/7i2vEYb+t6QQOWwwLbEts
9Z7SK3HMtoPX+jF4E1/RaxQUERDhvm2OVYRArDPd2xk9lPaBWGglXQnnjYu6nFmM
Bfqii6EVfGZdjLZKKFUxuTP84qIljanuLUT/0z3VtqjbGxnGRzfvcOyXpfou6sfg
HrOJAqOxqiaGIyrDrAEOo2hpxJEZQgsOf1RASE548xMak92IWpM0IGlqM7y6qPcE
XF9v+0rBF0qkX130m6kcDRcng9NyhtfuVjdBSLNxbdSUXeMMZ+KUufKAYBHr/LFi
i+Qc6V9D8nTPO/RQRTzckZjkfgsEz+CjZpQb49+qnMl7GLZSbdQMq61wY6Wxyv90
qoObp06nPndZuChkWUV1LdHnjIke7rMChJiRosONAMIeHUUIJfa5HOnF2uuQ/i1J
vtG1LySlBL3TPfZDfBqa9n+Tt4mdgVIpijVZX4g3Aimz5q9QnTKIzdEpgGVqgDKM
JfrWrCwKELpxsKZlWoBKJfXGbYcdQFBLpODi49K7qhIzPfvJsqGAhprGvbpRlmK0
TgQ7CEeZfwCerwqP1YYxoQaVeJ4pZUZY6adQc+cOea5UUpddkV9wc4A+oq2amEXn
kimZbLN0RKu6uVaCLlROWFfbLudBlHN+bv9JChDqyQlHBlywKMAmiWzixzFEa7ne
Rdx7Hry1xp1CPCExyLaHVX8pTJ2WuEstGicoVmdBfAHKZjCC1FuHUU9AAeewABEi
bZlft+V3Nx/7gsELjU4WmBUgjcFkCu6Gl2H4VbjaIzj00z0XQRPvQmXeBF9bWvNj
fSLKtOifxf3hcmusLk6ezYKTb8LncBNO0FktuJmZEq1ODLLW+xvDln51gNfwWS2r
DR6KWSyN4fKIebSCGMjCDErvSEbnSAmmE+6UL6SyBYJ6Erqcq/7P5lH7Bqmj4cjO
TEXYMq3alpeb12gmGTJimKpCHdP10/IIGJpf/lWNEpE68EKqBCevm9b90T08LTEr
xYNaEYsFscs0LI+WFxzADLro7V3bNdnGjG2VChMzaA/xv8gKK6drRmJBBBeflbba
o+MDhPzUDjxl6mxN9nDBJV+1K3lfzyMTifv7jN+yROVncHX/EDkazE7D29G7Enre
huxMKdomhLQzOyWIhE/tuilXMFFtfHwp308hyHBoGUKK+lEjRqLfX0/TbduD9b8U
WX0kGfzfBRRCPyIejfzOOrC8+PVf8OJrb2LUYT+jf2x2qVPNiHy+q66fuGndrXJ1
CVuTilrffcuG1jtnql4QXRwYasPLU5RrXdKgs17vJ7qsaz1BWjSWmFolYZ/9b/IN
0U1M1OvBrynNbXdSUye3ACfX+sbfADmruCwdpdwg1Yk6BAAv0//yeSFkLKNxijiY
ifpRcK21wZBr8segz+ImMW8sMcgLgyMVKPb0bDCvSm3RPKwCHiTi8WrwtX5dotLW
fOYy41FpqErMf7Z/R/6vbPrGNIKcwjW2QQ7KY4R+Hn8Kp92prcocNAtxs8FZK3y6
vJAQZL0Tp1BESFwHey8fyNVvVT1zw2d63PPAsitggJg8ElNdCpsBnsyumz9JUfTR
vKn06MVbwQiixhSkrrEnurfv66sMlTiuScudK4+Bh79dPZIhBgvY/bjoZD7Pne+D
flB+hm/vAkyx9uL1HnW5wsDqGEAsYWRfO1TLAB6+odNDenpGPuoUpVCNmt48yd0R
0Bnw4K/iOAkxG6J9Z6aSS74NTJo9w8j3+v6/6jfFIdJmdBkS6foEJmoDIvtUzPPr
tA2PQ4jtRmbYcun+VM/Vj3zKcKOau1mkFM1ukuomhlSqReh0mrmhzVq8rpE6L30K
8wJkpZDjH61M9ZjbfU+qgOnoB7qaaof8Iq5VmoHlrUcN/d5GnOWD+Azk7yHLbSzP
87K8DQb6l5gQ67S40UeR6I+2jyKxdYgF3PglwA5sQqVhAmfi2t1afg5f+CpFZBjB
WK4uZ60KtQfWi1+anVbhmtnBed1IhNz1RKm+BoeG3ApCRuOUCLZ59clypRRoXb6R
XIvHVHQdgrS3sySu/sIlGDJqBDqsIZHy9nwjeUwvHS//v8FyVxR3ZItRyrd4h544
adG4SahGUAAfXApAmxjxoiTFMOt+WHvCA//6mkCzCgj2W3wJ80mJVN8OXIG2mZzr
aO0pVdI8v7zmxLrNe7tnKEUHpaPl7LJGrHIZK55ltCkn+35ZhvqdDl/XfB4Q4k3H
TznJxMhxG89mwKy9YDvC8LWbHJRQ1UlopJXuWWFMHuXdFE2hTwLIUDisYDKRmQ0G
GZ1HOjBMGCtcqAcg3k/VdQdzvc4DM57If4TdxNw99SRSmhIGYy+sZ3pqRF2HbJJO
QM0bGZfp4KVMl4/5xT0N3btAXgUv23rdk04qDyvwLEj0dOvN/wN+0pZhD+Wf7Iyy
CKMyP2QjkpdA96ibmUtGNdC3gxMpHPYq75HPVStEze/XC0gW0bzcx1J6rO4fBFdB
AmAKZ0bUeXvRJmbTZmYRh6LowUEHpDCOPWO9u4NJGnJ/OzKyBy3YQqwbu9FpwcRN
guadVfYP4sSIN71o80MiyZBxK0nvGTsaioO0U72yHQ697RGcQCBQG71qLD/SFiVD
ZEdfeYZAF7aWiHD5RbsvS9QFBBA7qDhrAINGTULvGFWeVJUNyt9RrD5Zh2oncCH4
SPXpxIcOQKyK9gLk+m/pDX7DvH8a7tJNKjnu/NbdQT8z8hCqsJngejNTXbNTuP4N
Lw04tjspns/rUd7iKGjatptjpiQCOCBhw/AWjLPJoTEOW4UavTduhRTxDdW1L1he
BbuMOzidej4MzI61qOMHNRrj7N2htjP0j1aQ4egmSTK+KO+n50VZNXq1gVV7KHvB
mpfAkALMb7J1qWvQtXcG9GrGLgoHDQ4+z3nxPtzCzDSF83avcAWNLdFYHRZfH11s
67chzZ6syej/sPU/WgfcD9vpLkeV1RsihbOSa9gcgJEtKtDc4O7WWkbJikyZ2YZI
qFYhLE1FUsdXLlj9Tm87dEbjG254vrnX4TpuDiIQdlKCAqM8CfUlqc+OK4zQc6yj
EVOcPy9k7ZdWky50+kQIlKmU3tvbLb0g1RITrNIDisuY5N+zvLCCQHlH4Q/Vaeby
+U38JhJ0ygnVg3GNUdkfIXWdY9pBDGab5He7GpSwJa5uYeLyvJN7U9/4GjPScxjj
j2rBMJKutJgROeedZ2vfdOZyWSeuqOCGvTImbRp6CpaUcklNdC1XgbzyY7lVtBX6
smmTj6BtnDc1TXVeYVjDo3v+xv6Q1MlQhm1Y+hcDR4DHHk4HMuPuFaX19AP38xMQ
bHSmRpjmkJc3knPpCYOu3mEAZKN7v2XjoluhwctOBXoo53wlsHZbvjMohBdToLRG
e1Wx3lC+bSA2B4DClr1LneBz8HXW+OF4IgwAqNiu6kaoHXzo44Cz9rvl7LmB8ZQn
VHbQ0pulLjM0eDBHaVMwxbdxADUFCOTcDA8q+yNHJ3zJ2AEp9E4qZPO6RiyKqjAF
9TY/5ZuCPaB6a2Hu9xY2cB5XPAwBfzTLSi5mECc/G/PaM2FfGyBFeVC8wzdRGQ8K
NuxGxfMLqfwqMngh3nzc79DrJ/gu09MB5U3yMw8Wl1ty7joangWbmvVlKMBh0Tek
A/2VtjTPNcZ93G0XJk9IucNy217Cf39+qKsXlVyQmrHwyoBczEJ+ggvlwc/KHBEt
/cs1s0qA7rPy3Lwp8ZCq2ZW5HNMYXvTbxJrM31B4EGTQZ0B8AdhwWbqx+GnES0RG
L4QySrrsXcVDeU9ZsydWxwR1dHxJxdA6GzLz0GcLaQxfz5j+843BsJxuJ9bBNItY
FkyU6Ghj+S7+5EQOY6VnQdplHQOTqhTTgtV2V3oArS/53hmztQ4cAerG2W8wTCyP
HXeYnbeY66Mp1QfwkjOrHtIhUCbivJhL8SUOLprmW4x55fG92oOw3LDt2c9lCu7P
MGQZyY8jn+sVzKydRtJKwYQWoJFIaJuGywVNofDWVvn5oKRmoUsdcbi/3/XziuXs
YpNS9RsCVvdCPgCylDiQYCL2hUSS1dntsdQzRsoxXSYD41Vc/V0C78j+TrK+MAaJ
Dw1nWaBxnPZ9jhnMX0p+NV/RytTZO1AWCwC0cWxxU2qcdlsbcpcmC8reP8K/CBPS
TNQcQPDoTcdX68YOvfKxbWjKvyMvqQWlq60EfQcotbEWfR1XwkhoF3lz2rSDPFSE
gE2ZtPxfEKUTcmyk8SN+lig8q9h4Mhxu6w+b9kP5LXke0rXiMI99cqBc0GK8YZx7
BvB3bo5jq3Xgxg4X+51pZYJ50Ch4TMRTPBgveQwiXePELySjyFSIBnBTm9EDiUCC
J0vZy4QeIqWWbS94z/S4G/orihMVgEPmvi2JmQfN43ruwVHt/zf6wId93rj2tCr2
4FSbGfbKZC2KccG2B5ORhj9mb+aaeCAcpi4d4fdPpVIcAp99xzblqQ6TceRFu5vU
dMyaz3PgKna8K2q4ASSlBMkmpfnD9CtXteTLEJiUryQL/Xyx6WRI59RtHxhOcCIE
5uNC+NETW/cjLE07mlA2aOoPykmZvFippb516G+6MXrz+lkwqIQTgm+pYrfk1dZB
ga2ffYJulndI1f5pg8J+GTigmF46fEWgMQ9rFBetRBBhC/rwjLEfPP192md+4KL+
Zv26PrFCTntwj3LgT18wBtYXppXm9JQJ5zMJg8HmdgynpZ2CXRIp+V8rlOhs2m/N
+uUqQ3LfIjoyO/fqTkBecqEml1yRXnHhILsKcBZ85PGb321bfyhXGwODahyEjezs
PJzeur6+rWJaN2UJD/ZBhP7v/cKzvnUxoI/qaF3Pn5Urq2AHQZ+gJPwu011fGOoq
wputOIj3uWvSnAJT33tQT/bXjYK1K/HTBpiV81jurHaxKKpfo4KX+ppJ+OOdAj8q
mnWw1WQKNRJhVJjU7LE+DkfkFKfMGzwCGnwRJ5x3wpX3NsEDQvtZjUeL0KkewkVK
WoFyehcwNmM6FlESXik99t1dczLgVSaUiR99ZRpHigZhcVbvInhgyQE0h8oBPiMn
3BlINt+rcUxqnWVPT+6vXG3SrIMTv9qve8fV1pZeINJXDJEVun/kbp7c3gNq6JZ2
7wt0RQKk3a6Ca+byDAWAISU/SRX+JFUM/bxzhtOJ3+4QN2gihQZZuKY3XRCzaqhr
eU0Ql+bcn0gEvUspi395rkfI72BUwERtlMRECjaBqPWIGcwk5jEmO+SGvgLIGXQW
xnr8HrW5xzGTeEORCrM5J/1Eny28fVCEORU439koS9wm584XLxIaE08ZoxoJgH5V
2r/u7mwYx9KP6wFOjYHjfy/W0tLiC+k2PrjtNbFxQJkq3fBg3YjTiZzZuo9ULMXj
Qm174zsuJ6wm98AXDI8Xr6wPjytNF1RJ2jlZglG07dkRzH+xflwmXXf/mnCjyJtR
Z9nAJzstlOVzLg0WGvFsmi3W/Q2yAAzgELZkALOrjTZThpkGzFmuJM7fp/sdk/oK
xQHkWbfM/g9nwUc3TOwXPfusEeqTcW0YgHaUswNlnW/JrT3Lf9au0w3l3ewmo2iK
tfbubnKRQ/LO45caoPuGHDrhd2aMN5Sa2tgYGB3kJiWPapfsvlef1LJZ4fiVq8CX
ILVG7LOsHnDP5Rl8WloerTD2WgRll9ClSIpHD3EGK8HWrcUaj8WnaTn3lUhpLmGf
65DsqkHh0wR1YvRNT1Fg9EDm7jjBUNjZyALB0L3bm3Oo4sJBlV/myaKaXXo2XSht
KbODhJAr7+4W6v+xU0BFED2P1AmldMhhC/gPVQ9mw+U+5hJqCYkpANp8gzoxeJ9G
lgFBfZdO8znRhAa9tUwK7XvAQDTe+kNOKr86m/qZnC0sWxxhKyKpWMJ86/XEOIAQ
pZzvKzh0KuPVonLzH5E7Vl12YcfsqRcMmZjQ0zaPJU5e/B2KeWyKJ2BSxdFRMJzq
2HXBRCUOlvMcilNR95Oo6x5KHSFtB8+skMs8P4PwRTBI0tUAe2uL39wfgWtUwCSU
o7K/EVxUnXHUX+28oEw/A3KuGvH62A18FenFnzR/eXqLwte29Xcu/MDZZUSUMkAg
cqtkK2hKOebsZf4oVcb9ZxJwzRel7J3lnQ6HD9En2Xmpu/p4ELfsdLZvostKyiK7
c/koFSqSnznt04K87q4sFcQLDaLkLvY55nf+xLMiogCeeps7YKwG63pNY7tWMaaK
yKeB0vGYUykIPjFCqxpGmC1t91N7uHmuCAGh4vk7hnGxaRED99o3a3U8KnB49hIG
oEDRezfPlndjC3ddIXPFGfyUq8B11v8MNEEUOCBssWZYdYNXdh86gJTfHYFZKb/7
sqxTddn+0UO8Jt+BWtiWmCmR0pmfgrLxrdDbbnY/JxP7/elCDaJY2quk+lKdJEUk
RraFnSZBiCf04dLHfFtpSj530g4B6VCIS+3sjKlyaY+K2HjLmUutenSRsCaL3cEg
oUjDss4ba9zFlCsUkQ7DPbMHo15gDxrJ77G5wm2EFbB2M6YbxsfUwQShIerhnxYJ
wkWnguFpzJ0bnWTdx9oVpZjH5MItq4wTgHd56Ehhgbr9SklHBYQBukR6ad7YQK41
IOIdKoVGmLiqvWgmS+8F+LG8cN0jVnoJW5iFlL0sVOLbVLmDTOuIZO2BI/b9FEAc
Qj1682WTTYI1rXa1uCODOIsy8mN50HfpVvPXhjpLsZ3t4I8QJ2tDzdMY6/D0ruJl
nVWjWIXdPFoYBJPuapr+mMjXoi+ZlVeGTGzWNLdm0+NelIEoSfq1l5csUje7zRMJ
vbdM1XyMFdke4uiHmhTBqABPxOy8apZobbohU2AxUcphC//TjfR09t7oGEV660ja
mL5shi3+LgBkiPx8MLYCtjKQ/cENCoZv7GGlkyOOqI3hKM0LRPrLu4l5zUXRyhBn
NDMqRNfv1tl/4b5073sDWGvI67WN2DnoQmzOJp87Riv4D4bMPyqiSr5QWbquXY0h
E8EY/w2AMd3onvRqwF7RDQmV+3d2RKMS//QFvmUnzJY9D72Uc2DUCONg6hR9Glls
XHowruXW/JbmCBTMlrOH263c+sWVNPOxy8sJY3qFsHWTiFi62A68qQTa/1xees3l
3ZGUejuFQj84DFbIs5fYimShyylr3wF4shig03u0S9ZWiNWIBf7c30bBEdJBuME1
3xZiDiMq4WzmBjtdoW73nh3sdrS7p+V20/UFWODMatDkyyXziO/XfrfvNZI8klLB
Ejh6Yx7EMAE1DXSFw7lxnGSKhtEHb1EqTuiP4D3puJgCvhJctEdkyb2Nw7laJnxT
MhE9ID4ssIRNc2XJKpsPw9O7speXXWvP5dEJ6S8BTvTMlr76SSp2INdmsuN4Y0F6
fwwy5yK1JYwBdo/oBat7jJS7mg/dxnrzR/4ZYRz3FFRa3Fnlg3ZVEociCdVZXQyx
hGtsAM7ABDTcorS4F+9atyRJ3GJvi6ofCDuaw8DLWdfTSVtJGZotgSP5m7NWhrmP
SYZsR7kJCaUYeOjawykpmddHydpl8bRLS+CsWO10BgW1EY5lHkPC1DsDj0OywWqm
DWkvOoZ1Jxsnud3CDD/JbJJbn1d7XQZxD3Yf/PrY5zBu5xr2GEs1qJVunZdHS3Nu
Lt3pES6r/Zn3mxCoDWznUIyB7llyWORm5oTpOpze0IROS7iPkQSVb3+/daXhECmx
3tKnhLyvUZEtx1MW1SQRdMXQ8JvD7F1YT+aETWdcPy8DWka2ezrovjX4IvDV4x5U
lXhs9+7jamd5h0m6tBOZZ/F3zI2jAaUwSOwPRr9xLwaeE8iDQP+zb3XTufE/+tUH
KOOGNh88X1ExRseDbQPp5RldOTtZWACbY9oNJYMydG8k2/B9fcLOId6AmOB67ohG
VX/YRZeHDhKGxjUkFQ5exxtpEQ2cK3T7i2IFrC6tbbB0KPAu41mNG5t4HpPsfmze
Hj91yODh873YICYQkfGRKpRbonKkm08d/8KL5SUilSupUhUeovwjC24pXqFirQox
RSIwa0Nuxhk29pV/LKvquQR4zwxJ0XdID6TNPnDgn+ym6vUT9Dl015PcveT6VxQq
IaEQuNXeHaxkumILBiX7NBa/0F1JruaJu/isv5VwViVic4sCxAGgieh5Laqo9JyM
tMJEE4kiJ5uesKPjdgdQ48uKJ2NPxVd0L7UQk4F6wNsEcTzNzjJwkYWVUlqQj2Tu
na0UdZzaLIpVFEIS4di530KqXZUAVEvUKOYaTotyjjF9H5BtvsdZevJqZqq9m8Jh
Pv/2obFOmZ3gBP8S4tyvMGw/uTthjUTfwTbqqiR68bKrMK/Y2rDyeGXX6erH8eR3
ZiWte4UcNm3QE0s4R7de/a07LJ2Otsl202Xet3+/Hmd/T7iaP2JyvOPGu6g7WcEr
/i2g5tfzUNz2OXDqo5wEx6LBHJAOwDTEp9jwmnexBcKxVybzYwDdyTCCw3ds1KLf
R5Ar16/EDOeM47wqzYVPR0Qh4olgkzoLhpFv/ueWippA7AVzJ1g9OGmA1ObYDWxP
oqenFxqQakxg9pRTg7/dKYLGrq/2eIheojeAPU0Tsm91qgTaTcZneiTsf/E0jU03
PJqV+Ssr7tGdhHy8Rv4/3vSm5AFN6yNSGl4M7RcfJE37EgH+D9rUt8AtJBRpxHHd
xZGUQ4MPY5lu0b9qClY0fMnH0lQzmll/pPL1eUZ1PYneAGbfBBz6HseZbA95rG43
3QbE0yS24OCHkh4pI97IcXFiXMqM1459AjAIiBzbwg7BeJ+m+aRwFlfy/TjsxU+v
Yp8muILdowUm/s5Fyh9Xkg5dZxOF/jHkKn9E3Y8sCRxGGdbhsUNRw7f1l+LwY8MS
Qfe8x4dswFBpjiog9i+40yyp1RrSOmGdvE0Ip/ubD94irMvMubeX07b8OS+XXV7Y
DwpD26l8G7OBZImi8mY2IdQ5a9SG2n2t/k4jVGASmEHw/f+z+Vr2+zEt+nhg2FQj
vUASbsyYS/SOejyJxX8ymRLjWApIZc7FmUSD/7npkx3S2uJQ+45U48/gCxRSTqkA
gMoXhyzuxC3ilJ6qJL4UpN+y5pPtJmKn0oZpuHJseLYaoaFPWFl/q7MQ44BXwXXf
SiQ73zqz/KLUG0ZoSrXUusGXUNswbbRUi8ut5qC2Vb0TfPS8KbVxu7J6E8P/6i5v
I/aJGLFsvAD3f30pGRQkBFWN8wRqxCvCWLkPpxnFxuD9aV4C4NaClB1eLHztksjD
+gIBEtMboy2WO1IN/h4IBSEBBm1AqO1FHTlKhKO3YOHskWK+hLDqUA1zGv8tCEP2
s4FO7RhykObSq3DXNaxkI3bQSs7bwyFuQZoCfMXdDICN8vAAdUuDhDITWjyxU8iJ
5mAQ0oYfSpJ7eX07dvLU5Vqvi63cMs9Zw0cMp2gGlVaLoyb55I3gnbc8pGRftXf+
kw3yE8FPzTLjUuAUJpr4iJuWOHNhiR7tPlDfRF5LamhtMh5heQ5sAanEg4qaszMF
YbGW8/PclR6X4jMbYeYnV5shJvvrcfeHLyhlXv/999VPNal10nuboUgYY6l9BdTa
Fi0ufcQ/yAbAFA2uYdRoGuMmptXXIPqudDV169APACB1xVz8pA5R2F/X+qCkFVbO
ZH+GJwwuYBma5w9vWaJMxQ5acxpKN2BePhAVSlcilmrOdFbPIIbWQZLc8oVIhItS
EjsriG1D6D6Ccx8yFoKEiYRfExtVxaBt2hg6wiyojtH7PNvhJ5ris0lo3wekU7Pl
5OwJ4e2ZE2eMzolw4GJLH9bpzu6I7/WO7umUPxqC5qmibCR7JD62zdWIiNfReaRQ
fNImxZmCXF2x/UOC851l1njdqN8njVD8zVdeDtVuzR5WgHgw2qLBOa/SVBtxilkU
ZWnCch/IfNxytXrXfRUa/s9n3mLREjA7azL4CkQnVkkb3jBg6yeuaJ96PktP6QTb
ByoalfEtw3xdRzAcFtLPnWBki0qFXOIKLC6EhfKp32hfsXjbPbjVP7vJpX+KEiJm
aIhgQejlH32iJ6m5hOkaeRR3H1tELjA+632v5mw5T46Io4s9vvuz5gbbWdoKhKPg
+L+Lai+Kw9RJ6zNFmN5lDDvuwptGNpy6Wga8BdEmipTwl/QFNN7IdMBL90T2GRgI
LYD1CrGolPqDlDi84KLOAaHjfbzXJxmjqrJCQAJZEzpzSQNWgRkevdbhxE8uzqEi
39ecg6/8h18g6j46L09T/ldVdI0QOa4MJa3SqIvfuDZU144Jwss+/4DomuQvNewA
+AbN4GaO2zz2YwJhhYGp/RKjtj7ydPtchyzhCPOopwqwTlLPi/4wufulspqrMEAr
paeK4u0cbj2iOt0YIEuc86QUCk5pwulP+eNC0bn/L5kCMGPGpGyqqhI2nLho8s44
tyDgZiKjkhx44I2blt6BgPvEAXAD531vxwT1Nyiv5WkSbvsKJXmrv6ili7QcjJQd
e4YkyMUkqjnTADEIMFZNwqCQ9jsorvFuXBBVeQj4LkGKf8XpyBO9Q/4QsToSWooI
7w2Vgdq2NNBWg4OF8gH1MlQDcz+T/P6GzQbjrXXya5NHJFuM37jf8jhZJbu/hgKT
52s1+7YePsM4wsYq4lsf8aatc0niETjxlKOsOEk13EXGaXDnjQMmj9qefVKH1YUO
e5xGB2NMlRiUa9HWxVcq0IoXakLnuefMqA3wuiVNwnEh0v8YX4H7gHRDn72ikGv1
PS+9Qdwg2KYZt4jUuhPlViaaBIsF8+DhWSBERfUMB/hSezAZf6NLS05afF2Fx9VG
/ttcaV7LL30CnP0pZXWA3woTL7YXCHOIYJfSY1LWMsCPks4ei1WIawcG/Zpi7zKj
n8Mcd0rq7Hg+EX4X6DjEfO6jw/8IC6A5HL5Hg9znIDcQHH+iG/eXLWjVl28m6+Sj
lTK5xn12CrMzKRdiNr7XjvrcW2Y6G100JDLS8CPHBgGEeSu1blKbn+9mlfv+Eoid
sD75f+KsAUJWdrrOG5GvAhnhulO2A5WTmaWFxaFZ1BeJL0aFvkwLpYqdYNJousgq
UWABvzCjfbheacsyXCdzMUTU8VybPgd64mMYMljJsXb31tXmrsiVbiD6EFSuKXdO
BahqTLBrPqijj4O/acXFDU3whr3KD+UoNGv41y0hyE+Ltfv+bTn5K1TpYIgd5m57
DzaO4cRVKltPHrY8WsqmVQNJ6GlAtOz8J/g9XCnQ25pJulf4n8ocgoFI2gummVg3
LPZfTQedSaA9f53sz7rZgMs4WSwU10hEOlNKo/b3iilVn4OUCEZrO6Aym/8/g3lx
qy7xvhuhLa5sqjUyRxcVaRCOXXQQ5MzlP7EuPFFlfB6DSDha6Elgsqex9an4/4xj
q0Y9zvJvds7Jrlsqga+2bTdao05X7Qrj5hJG4kRdaOiFO9X7pXQ2YgURsmrhThCB
OK49CEnKnjnJUO8ZiSFPLND45wZ6NqBZYNok7Es3BmNfTrVLCGHS/WflZFdyGROT
lnqeruQRW8ZVkeB9B2A3d9w+htVkFLW7x3dJuER63AS8JfBHSbnvI7mtgc3j1ENf
0OC/K8no9eD2aul4kjdCsm6noMLgQf+YJsokzoyVU6ZvFHKLdMfeQ5FTylQsiCF+
zPwz0P+MNGY8VXFyv/8i0W+18IxC0I1kWb0We8Bl9IQCw7MPFBsXXxliaWEwQ1+9
KrywfQO98A4P0RWOHsywiT5Z1VqwkNidIDMbW8OlRgaZtJomZSQTXBN0RoL/BC+s
kAlHyYV7v6nk8OY+eb6Nz4spMj7vXjRK43uw2eL2/RBc/wUFqs2HDUb40ODTIUdC
HSZATBPrzNM4zxAsFue7TVcWMJvxJuveOR1r+AbtK0EPOVmRbLRbhCtN/JqPPejD
aRin+d/Ph4uHl7dLH4f4hpc8sAhD2hvgKF28yYj3Sr6Op9FZa8MZ63RCKjab0R/a
X3SH92efP7cW7+z5iQX+vmYArE4/K1TsopF6wSFjd5yVIjHVrUHETQ81Hc7kMmT1
scxOjkiAxSROoC1oqR0Rw20+slPPchh6BlsMcVoXZJsx4nMCgseaW4S1cNoCoFUP
h50klnEaTiylbLsgk9e3vdSFDGGRREZ4Ov8bTdYNKBFSwYff1xfdz+PUKF3dXrI/
5oGydbHWtoXOMgoI4h2P3xXXVYI7JK/PtRkY5u+Jo7kVMZqmTePL9Kjc0AALid7u
PY92vHINkNdDcC/oBKYmeUZtoFzsGZElcD8LYfP06Q+WYLcSW1iuEyyDwXMSNDD8
Fy6wE9Q85qRaNrU3V7jZyTucSbBWvgLL5FoCyK1teeWYrXHLOr+Bi5r6Ef/WlJBv
4n7Rwso8E9C5hWngQLr5CyHmuv0z6EnETA6PAaSsdc8UHYLmkeK30LHkLUSnA7uG
HZPFMjQ3MSZs3U94jRj8ij3Y9Lbw9q7yvJYafUURQmGK99t4f2wEWVECpBS2kbgf
9HvnCDQwb5IZi6TFZjpgVwEhlJUiGFkgcJjH25NFtAhMYJ5fMQttrspkpFukDrFc
1PcY3vHvnOx43d8lib81W2M8q68FnIwwXZ+thJ9ee1Y3Q3jEw+U+Hf7wo2vXJgTk
6QP9gHrMP67WujSP3pcmkAeIFR7dxE8yvSan7iG0PGA2dkm0naVoBeRyMuNT+hn3
OLAt98QxvizFpECOep/1X/YMkl2umzAJEr7u4PVOS4wUrpX6zjZT0M5ghCeN1CRR
2T1eIji8xQJiHGIboeseu+rYPnd9FgfISgiSfCNicE/vuBLdlZ4/bAhw7Y2QncEr
/8quzmO/MrSSgQGG6VVvad5W+hxonNsi78ISYI5G54BYZ8+oDIoNd2w3MbEGLqbt
I02klPBgGIN8V5iYo133VVZM4c5RO9SHkpUPBqZ8Fp0igCzYJaKoBKkgvxuDjPhP
2FljOb0LtZ046XBpeu4R4XIVcDr2kuD2In0X1pTffIyRH/9r/xz7+s0aPZqF5NzT
9YnNyzGe/8DLD8u9JbCXZzcPRKHG0Jv7b7zWQUEodFllz+dDDSVmVUiQVV2vrJ/R
mxknmSRn9lh/OlZf38/whWlSAvfQBuOTdwazRpYJvPl8erGwb34nUKtnWjKQAZfH
punmg3Vviy5M4I1YqbFfOzJLWl64pmDo/U7ZcvKPkn1Gk/zYl91b4Kh6PiH8ywoi
R1+SAHs4h+flOQdys8pKl4hy95T2Gdd91znLtQUzirCtCopZbZXfIgyByMjDxB6G
/k/H87P1mTsQDx0heGFEdS2IU2obqIN++uFP7kyKgAa72G0MFi52f4eUbfADMGbx
SFzSNqBzqSSXW3dey12qXiGZjoEU0K6Z0dzzjyLajiVcx9VlLVPX/g8FPd3VKQwr
iqNDoU6sxLx9bajxALnvIWYIBVnONX+EisuR9QmfLqoHEEvwgWbzBZn0DmWVXXJa
2J2zg59j0Lo/PSHAtUp5MRiytvt4krGw/fPthTtdaTrxjIDmfnaLuevCiW+xmvpJ
63gUCsLFkCy2qYb0zP2/7qZe89TpgIN/n3+LAubVwllLBtFpLFn7aI6EaP9kCIkP
zU7OBe0INIo46PBF4oV+OOsEeIVfJgR6R3TcSrF1sKnTN2JBtyC2iVeNEYCGd4S/
XHlr2919SBfkU/LqdRk7S3Upd1aQEEbBP8xSyOsbA9uq8x+CgTxs1dX0TKIGXFzM
6AUMliXXNQcI2OIPVsoyCPAGLR/oR+2DZaL/aw2/5f/iyuuF917wMvvG2E41bHZS
yMVAL7wPSFTa0P8WqtDmch6P+SYmtMXFD23lLJqrcbqH3sigyzL+o5eqK+CNRRkV
y27+7O5kNvD9MU6pPRtfwF6ktdOTgG+bubrHog5ccsRDMMZEK8lXiI3Z3VoZ+xIu
Bps9KykI1jyTk2R8jUr6H+Z//IwcfvLdgIVs/x+p7jZggl3VS15JuuWAZV0WNDkJ
DtN1zYFfTaDEeORSzJg9gmj5E0wRjCMSvS1gP77MBlSAGh/tX9RSnhArWYioZIhR
cnxv9JT4Pz5ukM1UJ5aT+mEIE+k/tj9cgEKy3U2/jwyA1sZD/SpKQSV+cpDGakEI
A8LSD63s39zR4QQbIPFJz0LH20requiuxeUVCrnzY5KiotazTGe40jCb6kJWXwt1
aq3lSGGUoOmr6aWZrRj16fQmMu9wMrHDszO7GSBycQ5u4Euz4gVtUEV6HhSHVQRa
1TKsQcL/88s+afY99cLW2mxbUQrDMSI+B4YB1fjhZUIawNFxOLI0+C9GF/lJj8eX
K9q63cJpJD80ZvEzVp1OZNnrbROYA5I5IqGw8Cs78uk9bNiuYi7/WOdwEndh3vm+
RDiqOWR/oCdGGiTHJLUMPjfeDbvYB3UUkU7vU8oRq/6W7PxTnWSHtEIsewBN02Vu
NdcKZUItN0PD37zI4U4DOdyHnHPau/WCuwDUN9QMIt9LzcW2kYMoeEragdz+HVi2
kpxjtPAxV49lQiTH9M/XXGT/aOJMOrSR3zcRM0iFhGxyWOcdrhCBcD1Dz/oQitso
febEZLP9x0tNv/ViEZxsOpX1RZGYN2zggUrlFv9G1D+wEPLZFVHF0+r6ezu3tE3F
wbNVWquEkbD5xF1S2j6Szxq+0SYO08nLod4WBeVN2KZIzzZXcnZVxV+urUX0QKF2
SeIUCH+O3rYV98D1ZfWqyJwtsO72BfHmIosDlHjPtoTK8d1MCZ6noJjzCYDnygF6
z6VkAwlwM8kMQYMfnMnbFRQU2Cw4cU1X8gcbc77BeOfCqxWks/pWUN67ExVEovTB
UvyBFA3u9ccSNngUrPMAMnw51Y7kbYn5s8e3WOPZUJyPSNF3uvf/Ay3/0PCAIMrV
X/Kjkiaj0GujsFi8UdTvj2I9LEz6egTCjBxtfs3qgADsDKBw1uMWkgvGiunQi80j
WuSDDIw/Cgx+76S5U4IUXFsqkn6L9YCsU8PRebfNVyu9ETPBONUscI2ZHDAgvASQ
ljMGyAlOCuQIikThaCFOiT6ZOPJlN6YBLAYwEw9crpyeo3ToTqki14pfOpmewQGR
3adZlkjGUpU4GPxH876t+g2Em2fL71QGll4oBVy5KFP7uxf07LJldZF39xug5wUm
kaHF8x+ENYKvaf3ngp8nl1ycBARdCx5wpaKeMMObOgun3IvgJ5UGy6G6aCXxNJG/
srxM6qVRuRgaHK7lJBcQrnptAmmCuvQGh9fcXXzvEK/TcQS5QWeMb7D67t0Mjcwc
V4ZKWGtc8mxPO3LCNJX/M64iFNFr1IlM29rHDlZa9nzURxoxRjhqLWSTPB77U2Wu
9234AIo80TjJkmMBNMqnHpj5vHHfCKROL6gWtKkSlMblNMns1W8urrR+PiVkhf1C
mEw0WoHSnAdv9g6oTDamySg1tAMKkR49QK40POCvL6Be9BTdHVggNIFHIMfV4Im+
Q1Iiiq68N/qTBZtPhQzsDY6poKkONaCr4vObOjFDFcOYiNQB4to++XlZEvTzCtZc
66Mm7UN26Pov3kDL27sOUyT7pgtzNuEV/K5g63II/6rMoRsV+ZI67jd2yFAhrXV4
58JeJIe8D5KQb/GWWrQk5ea3JGSsl9MuDasP2OPInr+4nUmkxNnJvfb0GtSzCY6M
qxk58lYlyzwlVc9pxXgPGBwxW0YEmtG9qd+RT3FcYA4dU70/fW9FObka9owEEFhn
QDByGgWCf8kOjqZR2JYgJ5o+Nqd8T866RvNAWMGpvLc7QUhW1Nh0pf/pRoY8wsXw
MmpS3G38G/EIKBmkj7xLpnltyHkHZDH5mHs1T8saP1khMuPMK8oSr/Qhk6r1ywS4
UAtS0SDGuko/EKuPdetLabmp+30LZ24LtxVKLyo9+ydim2wfwF+r1sS0wPl/iQt1
VNKuGUPf0ccg/xXVx9oy8237RDdJM/z4E9NvfW4cbqQESzlecALPQw0gKsqpamfp
+qwHQPPgEQWBRsfRoN4TbTA7XELeHW9n/BhT538agBQkP75vlyC2+gwo3K2UwPW2
EltS5EUy4QH6du+vJ1HJl01U40kBjpLUR9bno9tJM0HrrUUCT6wXUuloiSQI1njk
Lub+EmRW9pQZ5ezeACKdaUHW9Cn4im3wB9Nfg1n/vZm7i/5w0SU4F7sI3Td+yBm9
9n5MbDf6UMXZ8sR38KPqpuMhKiTCvoI0SO7QkciYxFPePP5Gt/uiNuP1e6retM33
J3xVBCQl0DifS/ixEZxuR+lR73H8+zAHHirGYueMVNQVUO0mpba7FLNQTNgZGj1z
B5KMXvHK6l4wOJlPcFx3exbgLCqh3qp/XJVD/7KOtkAJXP7EoCLZ4J+Yl8MTgDpL
/Nr4jdyqWKYfHV074/OvEDgSid1fXUEaC70aPBYZsoB5dxZmoUab5EFSzRyqjXiV
WcZRZwS68LPWGlMVcee+9JTptH9hIGwJxbyjVh4MLqKzDEDu03Bez+bZ1wEgfWBy
gFcxPXyHnNfVOHIuq7UiY8QhWCN+K22YXhaQJiC3ln+XZqJIQSRF68reDIiYgWJc
uhGxgkI858B9gQBK6pelOyGMGoYZQVnajeLZkGdomaSSxMAnTl3G/qW6d6BVUcHM
unr3U50TDKzhuBW/1fyUsYRA/GXboD56OkVRqvdBBaFVatsalGI/mEExYveqnJ3G
acA2XE1aIAR7VdHZDG5kjZK3sTrj8fEvvOAHN2G0d+phzJAgr1f0ECWwD5yZSo0P
hN5zLw/T+9KjrgXXgXO3DoyobhlycdQKm4lvjAt8OBv2VDsjU/YKU+aV86u5t010
Mvur7oYlQb2S+cBfpwhrUJdMF49lrsoUfE17h0OFJuAmwMN5Why9n6BXySZ0WdcC
l4evqDmr/9FovgH1agHKQIA57kCF4RHLfG92zSKmA8zyMpbv04sqGdoihW555Z1W
mM6X/ps/NefYhF+5JchLqTF2tdoZUCoZv4UR6v/ERaU/LRWKv3oPpbUix3fH4dBB
lyThpHuy+/SDwjS6wRSoZ7Xo3r0bljn35Yv0fSZuJBYnGI7zkmKUGAMSFk9fSPCg
9vf9+0+Y0JoxVS04QGiXmDaoey7QWpoiPD9a+SR2SCXZbAvCWrB3XWbJIycxEXxx
cTR3Iv78RJajZCaTLRRGhHx88f5srfMHt8HxiUj6bKAh3tbpCyVCHrasotCaTkdW
gQuxQDzCDPLoBaCVcCmsfbbrO1sFolrHIRi+4qdSxPa6i6ZU384PDnR9yJ6AJKIs
HrTWnutn5EGRcZOeuQrUGoA8XGl0LthtMR+lwZG8az5NKPZBF+IKWYCqoHBmPC47
EfUTnQB59q1bClYFIdfm75G8yBQTZbtLyMKdV04vKPd1yNW2hjs2b8tx0m/t3gtD
2hoOBhYy546UmydOFORfLVixpLA9rnbwUi5AIiAm25ecMIjrBUO0HzMdh743KBcq
O2jUHMp50SCe0fFmWt/RKYpoMXii6t+Re46sUeMONMWbdiF7KDakjAVb/7TL/HJ/
1TGZlY9K3vtxwuYB4iB3x9LT4pRoy+3FDPZeDXwEHd27w2ynhvGJb53bZGgjto1X
STt+w98dQjZE3Tdxd+LDZkT3znn02T6ofdpN9hJT4kaxF9fv9MHAFRhxCerVAyZD
oPVEDvFX7pS1qX7/duTlI8mWztz7H3QYRAPgWWa0QmRynpab5E9IXHKNGoWPRk/E
G1M0ItMIVoOCF2mhdk+SFImNTCwMJdZHAJN56N/dZFcUH55UJovjzqBVXt3YQufK
s07qfM9lWACOAybBPzORC758UKclsoPx6798a+G8TCNkn246NaFIrsDt988Cy6JL
zQCBcOM5e7fghJUtZO1Sq35NZTWLYPWU5nH1z94Yhv/WM5FebT8ou+GTNqe38exz
I29Sey9tL5uIRhBoyk2cImWIqReUV/HCDZ+YaTFDIWYXxNe5VF653jl/nYYA3/OO
5at2MOSvWFM2S/DXuciGYFnaBg2JQ3LwzxKEj6TIlFRt3/PUr3+91l/hQkKPqDer
F3K9/OAKUfu8vBOM/hOWJ6cHcVQ34ZM7hUIYJeufYyyRs6+cVG8y5I2GC85ykUsv
J1/3YNHEQomeAzfDYlBIIvdX2uy+S3L52n4X0R4MQFhTpLLGwrZeCTj4x0JbbDfc
Ee0TjIPPoE0K4SQNfLeVj24ZQn9qJB5Hbj7dNijkrVinio8A286TRw0fqGBp9ATH
z1g+EgJE/BoZBm1wLxjF0xpPlRBatDIjFgRhN3mFDxpZkWZMWUprfTIkf5zXP04i
ArDDnUYVkSSZS/oPach+QhEhd/OdFEyrUQF2WVGuiWfQScuxBZ2PrXdzKnZIsegu
dfCZ17yaoRY19B1cy/xsPhqiA+32mk582Hu70ytztkJXxcSeGasK8ZjLeDyXlZZ4
H27Y/FJ6wlN6ERS2QzYokv95JiaM58rSRQP0yu7mZIYJdCtDuyB49zgSZqkBUji6
MzGe0wOvXgzBhp48/xnI1PE/rhVCt+4/nLNLSsKbmXU1eHAyZpgquXccGlX7v8d2
YPog3VQsbXx7IzfQxTWPLxf/Q8knJNpwIruG+Sp00oMGLpGJEIdGCNohDkg9bpM7
/G/v09w/VXk1hptotqA1E6qT2RL60Eg/5z9wQl4yT5FKSHwhVzXWUfOgmUF3kiwm
pUt7TIdNZc8biMzOujeB7QBchKtPByv2EduOCTOjp3s68lZkGeTjONnDDJxAUfSV
blWeJlI/MQ0qT/GGbShhrNZFys5QmPZ47AS3KZaGoKYntQKeKgMTzEdygqV2Rsmk
yjhcsL3P8rcSKDOTELHrWwiBJKwC1RYdvLLYhIWjahLb1TdYIdNMOeQDuobM+jx2
SA+NMdqJHACbjlpLuUiU316Xzb3Eb0tqdaRbpfZUyoe1d+/SJinVJgyRNuWYXdnt
3NawUROxod14IlYNqBEUFCJfYv2JilM1oXkmQk0yYkRWOZ56HvdtLTC+pqaArwZ3
YG1mG7gDH3hdLxKhSheS15WkWMoB/IfqBCdh5om2DtWMfvAYaxhw5xo7sF3/7RcL
lfXajN1Cq3u+9KiFP7LUOoSjEd/DImoN4Zbsz9V7qXyYVZJ+uj8MB15ixidcPCE9
Jm8NF8Cr0u4FHpfnI7JlIPkmXrztm0xnEEPTd40fd3aNz7oAJ8pTF6yYRMzcL+TT
Fa99uHth04PoSFbdVWTB4Z7yiulpklgf3YRq9rXajMUDtCoIhgY4+FJv+AQkwfTp
IZ16/7a5FznqBjG4HT3TYpOZoZL46pnERQAXi0/IpjTpYVCBSDZLiyD5sUp5480m
gRVGytGf/dwYba205VFEj3KC61yR2CS9a2pbhcmNfkLi9gGHMBMCTiMxINqZimZ2
uJpm9EQaMCYm6tIiLunKnRD/Hdhc2+7zQuKQqZhUwknHDL/zVvOBUsctB/EqF76H
QMXL6FgUpfKQLXxnHL14kRd3rkE6gFTWr+eWGtJfIbSysFzQBnemCP9YL0GC/zKA
7mxczuRgKkst46l2L3wo9X+48ttnaHtbwopZYIixhusrHcrYxqnvo+B4HL6MWwHN
wSaEy8+yRZmtLmVc2k2ty9p+J1ZBZjRVlXhBUMtjmu0ls0VGMB29kXZda9ISdGJ5
zMjnv0m7SvGdnLGyeHCIK4AWFnV6aWf6EqWZGkRdkFvmkE+Wap/RvkqUnAEA9g7B
QfOgamUxzejC7g3MSaoHYy0sqddeFcUAQ2+q/bjmRgzoLv87h/2Rj6yGudHuRNw7
dEwcnEYjxkSsgNjvZMPr1UCJAFwrvREJp7DfPSKYbiFgD3j4fEI3Gqz6KQWQuOS5
79ReWXDraF2Xn+ZhQPwrRlZAWiSMZ/ZzTKHFq76FukkGBLyj+v2OlBEcokgg1kM6
wHA45MnooXG/ZJXMy2oWdP/KAdVhGQ1YoXOp662hggfwZqNMQ73Z2WrDo05dEh5/
o+BFiq4qi8X3lN+8ebeMhJ0pv9f0nXUZdhhlmfAlQxQL+hL5Amhi/fAsTzeUmdQt
3fFx7WRqKfvyDlgZi+GlKEiyGyQmQftykNozFDtZIBTjSWzqAbFp+TsCaVADc46a
r8EvuIU3/Pc02i4z3NH80FyL6Kh2pwizFwksOiSs3tlkUfT404uoKMx8Wjt+aOHa
Fln7cMQMazs694l3d8P7H7nksBRtc4yZ3Ah/Fy7AcYQzXJszOn4qcudGsZ9mB1x5
v/iPq6Z9LVL+sXsFdWE2CB0c9zHZtwyiKLLimwdp9QKKRRcyuaOXIBD3dxgIwfZN
tN/DHHGcg92TydFsBLtyKX25Yv2Dr02ypamZLgWd9cqsbAurBF2BLBt9oruXWPaz
2wR3m5pO8G0K5CdKZHhrQG+pQuS7j3gb9er1J36yBWgH5wdH1uU8Hc/b/2YVl02O
7z75zvrOKoHR0N3t84x8+9KpirkiAEEc9xDYD8AcR76rMl1bk1asqFS56XJF0ieP
GCWWZE+80vQDExe7vgFaLEwwdKsdicxVtQA2Vf3bhy+n3D99hqznJkTHBIltewnE
wSirUnYCsC86C/Y6r1NDriTvW6x09m/LNVdz73I5TvHX88GmhN8/C0kLDJ920VlP
1L1wES6ws8MV4rxxxmf0B8dCAqxjUwCe27jR76humeiJWC3eQNV87ecmp61LcBkk
kmhnOsUQG0aKMviT4UrjWHVMipLKuRmGxQkR+WeVJdSJuFR8zg1Ab0dAABT0Zj2f
/Hp32BW/MKHMex6w6gX+XYizLPrlimN9kFpEUrYmN3zhjFPlOhu6FCaS/JFl0YXx
jpPq4ubiuljw6cN5d0WWbZ03ISZ/VtU6MwkRENPNSyQlutmSdeGLnfRLzWpdEBtk
mXPLQ9TXyp2FU5Y7Ye141tiY53xxhIWniAxUGPxHQV7XIKWNI1hacj9r54AglV4Q
JnNR+XXXXgSf9lVovRAB0FsWcGsOAdtcbFpMbMlnOoF7AZpQTRrp5R4AB+bWchxg
jhhn7HpBoUTnWZ9bDva3nLTlTem+95AqUWwjHnMKD46BmQbBVavcJnl5hskYILti
iML88pTy7aSiy0DZ+TrjhrcIqkM/LYNayj61cy8Qc/M6PfyjH2j4NTQru2nWYruK
tPraQjYLAllWEYaOGpwrtwWaLObdfhawmvcA+HuldL2KZnz/+s0KhT3RW1o/9xYB
beSll6i58MTQ/Ly4yU82IdWAZN2K1pDE+U5GBbHpNR32JvbR6mCaXlKdqNtJtnji
h4fDCi3Ltv17MfhydEVLJJ5ZfATsB8l3STDcw2hK9u9suUMIIaPcXbfQPLl+oVj0
EqFY0VPcLI5nOw0W+RP+MSMUaRz28avaKikfMrodgqIyetixrM/X9ipZVzyxdvMD
Z8I+j9ocg9NeUwX9WsjmP+KAwkW8IAq3feaZASVPS8kvw5vSBL9r5cEB5mJadtVX
W2zCeR1bKB7EsH/51hS27bhRVNZyEbTYrB5oHbOnC4TrBTQis7Fs2vkl3v0sGLq7
rliK9JONza17hYGOlVZwL7eEDBehmKtnh1Sd5Vmzq1uYv2nWaUN8a1mo0vj524g9
Hji6PG+yVEoWrLbXQCFQqt+VkovK6lefDJ4ZafGArOAo8xv+MS6VMOtm9anRbZxh
TrKfeaJdUQ39LJBEHHZGJf1eod/T8lKj4iDKtc+NO5mhd5t7cYGdNej9L0T2sMaT
1MOiasNtftDlCdcBiaCL5a3/GGX5rpxo8nuTYkpt7evFeU43GN71/kgW7FoF07s4
QfRfr4c14S0fHv3Ogqdit48tMrqf3UohB2iZEorphmqXe/i4zSa2JRY0IOEc7pR9
4lw9tDKNG3mUyZBO8dFPqUj7Uq5XxRhyYAZvLcmdrdiTvM5QDeQj5B0GB726id28
HuoFYQ7uJuL/bRxCyt6J85AfEuTjHZGnF1DQ1Vfhfp5dCNeNVqXPTITtv+FLuxj6
eu6ZICxZosMdeEbi3i5HNfpkl7D2+nBzzTmEbajw7ydMfN+S9JbQi2eF3/Ko/1B1
MqkzXpRjAlodiWVv1oAKFpVNyYkgIFZXbz9pMDqOi44KswN0ai50rTI3Cq/ScTPP
AjcZZcMysSqAT+0f6XZESsrQ5I1rZlmMm8mMOIG7K7nICUzKnFoq2J4oBCVFOZjH
7y/BMWOAYmxpAzw+4/tsaoZO4V6B/Sx2y3vuYe9AV4WIIrjO35gVzXKQxau1qNic
FAtWgYXYYukEvaC8fXCXVER6Xya2BvLF2gh1JRk8hIaKppeuGdZyAU86ctj8BKYR
tCR+OarVnJJfEfZetdMNiqT68CcjCeKJSz/KbYIL0K0qPGqvMJ24rx4GPLN1NxNq
yZaOUM3PeyFQlesCQmgaW0ROrRu3nza1UG55IxeVjpUdhl9yNjuCPH6Qyqz/aPuM
ZA34auazZYbiZNwg/G40ZfPyWtfyN7gczdJJHygYbhzrbZBfGtY8QnG9bahMrQxG
/C6QAKId6W14inKdvYwCUXqzNyHrhkA5cWwU4NVL8i0IVFEiVZ3Tcu1LxA4fZrOC
1RN5AahXytRTOx+1LOPukMTMuhu54sLKbdW+GKZEIle+fSb9mrd0EgO1Jp7I6+wX
iC2ZbMt4RGYk/oQltpax1uLf+57z1e+MfXLvHLzG3J/pDbLUrOZ5TOHQ7ulBLMNK
btG+87UyR/0bOQ/mIO6alFp0pzkd5tkTJNSB88UhD7yZlyvSDO9euY17NvVOaLr4
S62RAPTCDYQycPDO4Htcpo+lQlWOSisV1UJdntoJDBRxsc85VhOxw3ur0RoEzxXN
S3WeGm7o5fdnp3HQ1Bx8ksryQ4hpCVdJrfYT886b5dbpQME9GXDmGFzpy4mENCQg
BSa1/z0AtDfWLAAMHBP38Jx+Oh1inMtzUQAFi7vnLxJxJvxJL5lwVc831DG8/9uP
O/hOYUZzauxwFNKkXSdLOBD/gflc3rYKczPd0L9P1WjGuer5ZA3oNd7QUHmmFlhH
opqhEoa5JMlv3zlmyIF5t1AZOqnsdWGF+O72RylDU8HQBNJoew5b5rlkrFA1bvVM
24oak+qnNJeid2Uos2N1LhVPNFRLYBMpv5kCo5ew2Zw45lSzvSvUnk5iYD+B6/Ua
Xp98sq6BwCSRx3s1VN2w9F3lj1NpITba0zZxQ11fqDQNVAb8elneoxpXbKIFrnkA
NyteZKZNZpQ98jT5z42d0eFtI1rmOcCsTSie3r8hcWicKbnPnfGSEkkT5bMUbP1Y
mN8BWiOj7pRPuxZJ2zVKQ2dAUyIRQ23UxnMyx6V6I8UWH8iHvaUuWQ372z7TCQkm
SggJhlUN60YPG0Xc0q2Z26/HVVkgyyEkYqjZo/J/CqRRW5rZgdpHhgP3GHPebJDA
V1pgm3K4Z4LObQSJwhKX+j7olvIXV9t+uMR+Y6lQJpWHqgywHYcctjeIxccqJrQD
bH7WmYYbq9sZGfJmsUyutipnX7ndvlRZuA47uIo6JeK5kw322cXpcYBzu9yoM+64
6sXC/xTreMe86PRlBX/LSjhfYROwGUaB++8Rdw8rcPhYslhiW0N9FFWffaGsDm1q
emHvJX55MVIc9ue7VjmdOou3CE92lvp/ttRku7kuPzh02fOSFdV9Iuc8sc2QaAAW
jRFEn+rMPZBZoQAMA94C7OAH4uvz6FiExVCjMj3Hg/lk890BurJttoW4t23/6XpK
liomSJLXrwP4vCO7ta9avJ5xLHKAbysnJhD87/n/r6VgzxQNxEyQZ7fM4QsoWTxy
kNhlyk5Slh1BaI+Kh28Wqg7vZyXV0eI1n3VtT9p4K/+U5jAE3hqnv9d09gUJqcYi
unmLeRgFr+tYoNFk+k1Nv6UrarNBO5ETOm3hUpNkX6ftYOHvQtvmio2qXjR2Su6F
jn/R0O0uF4n7ZtAAbxJkIulN6Oqozew5yTeLI37n3Rk9bm+ixMDWWzXZMMoiNdTL
RZEXmquBLhjyMEH8QGsuuRPNJVWkxTh4uO+wwi6PFgzmUxjXG048o/ZpLBDeKMQZ
ctoInN/BEvbRhb6Jo3Vw1q4dw54hD8ZQLYDoyaks94W0boJpFZ5MBJ6QHCvicE7S
qJCvs57WNkcUGa7T/4qTiTceX8iz98TS5cM1iaak+I05Oe82eNRRw0fyOrkvGo5l
/CT8zbzseNwEq9bMc0VV3E2g4mf+NoIYR8t8GkGBXMPetOrIHhRZ48adTJEJ7Ht1
aGIMd4UQoBqwBOiStuRhsTUDz6WU4xKWcckh3Zzge9JYino+jCmNSOW7XN08oPcF
Th+ZUQP68crT94oHQ1TFAT3ontSsVrX87TleQdjfppn2P44bgQLZaJU4j3VnTRoU
J7LE/lR8jFfpb1PuHFqLJ/dYJgo1SbS8uAota+Cbz3nl0ElSCMycHFU9jbUq4ZZq
gKjNzwDNYZLQhSNiB9CF1eA0e7i4kocsjDSk3Dcxsy5Inbq2tjjMuNwcGmZ9WyWZ
ni62x+/bPpWB1e/Ya8YtMnNGELItYK6CIk5gDMbFWZM5hG4tnDYajz1dScTQoFct
7bgS8AGj6DFFkJFhxAJXGlYAakQMtEIUwL1aShLWfGG3hRHfHz01T6XRr/hiwmpN
BjmwG2RRfBYAX9xJNtwPgSV5lgDpODOSeWjvEiSylMz4pPi7jMZZ/Six/s/nIgZI
LiA/O+ZxT+Uxz4Ghm5PRdt2mQLlaRHZCC+MCmSAI8c2zbFdN6++KNiWPDyz7z0or
vF8p2zMoZPN+2JIfMJ1UVnv6MRSK7fZUrcxIVi2Kw0KpMgrgFFts+Icvk62/1eBu
5WcratvTMd6dmUlmK8F6H26mC+O4VR79P9P0GwQE4p4akGrMW5nECG6sjp/4rGMI
LHmxr90mwK/UPdzz/vt43PoJQb+0XR0/JDictNFcu6IdawdxyMNteGTlU9Xq19K+
HS/a48PorokeA//HBCNBa06Dutjws3zcIJxVgufHBhX54eX0GvqOH6fzzd88i+8Y
j9OLaEamrhsxCo5/sJAyEaMOZIkRd5b8lix59TOAJdvTC7yAAPxXBdbE36VI2Ajg
NRAA+p5izcY2xbugkDirHqwJPG22Yr5XF/+SygOhlWtJ5La2Rzgr63GFA3NB+Ick
rHELvY0vDvQ/8+YXvQeUezjsR9hXp/mlx4eU4NIkklX0DGyfQaDARShQDPxMzqen
plbulsglqqXtwnLq8LffexcdP+N76H+0WAoHjFCL7tSZUueEF6lA9DJkO6TgLUFO
Jcnu2EbgP52dDB++yg/4YnHyuOL2AXpd5xUU3TREfn3HS6Z+c6codTI8XhwWYzNT
zRaZheq8YkrHpf1zwNsO0B4kSknSsrDlfW7bcxfv4baL3+C0rFx3cu0MGXBdONp+
m95hWjIc4PqcXLSUbGBrUEV1jQ5UfmM9DfsQ/1hRG97ecaSu3vV57sVuc9GN8KSs
Xx9ANgOcSYfhibTFQhU7ZzwzFIooAucFmlLKjlYgjz0SF//aD3VWxLqf/qr1SZS6
tyu5Tv/avQYVT5jr0E8+ZIOAnCtzFJNc12v54sXFpFkxq2CxVVWO9e3PyIsGaMHE
qbDxdsXUj8/Iif0UAk3RiLRQXtfmoz6kD6fiEeBwgxfUS2IzT5s70VDXqOIvUCVR
iTCoFSATr8Nh8NrfZJg82wyqImM/SUIIACuqbsTth10BEvwh5UTsjVfW277oaYGp
4i9eCmhFlcHzFHKeaIu8FqqxVQ0zrhoLCTGF4wPex0XBvVH8XKlG/v/lznu02Qwr
QiGJYC/vHSzUgMn9MHqRnDhsscX9w/s0t3/VU6CtcyRQCshF3QJWksk0uHgC34yt
ieuW9ceoQIeLVb2kf9QUdaPRCSC56UUa6II6BtN9fnm0tLhYOjje/vV+WRh7k6jD
fbAZlBSr3EAWzkBRc8gxhTpJERcnBby1aTGmz9EhYa5Gd6fyplglitIhwFHLxCug
zlo9OPcrgRYL0vlr88u7Yjmg1S2z9WYkSTw9JU5fIRc0fwREoXmep6Y1UQ1L5hlB
HcBer01XMouTQEXbiJbo2IpsLVia0eSiG7Rga30SHtCmggu8J3qnAOn3/m/7aTXa
1LoA7zKN/EBPzoyunLVkPgNo20e2Md1gWidYjHWrlB2LNVBf2lwOPlG+eMBDGFri
+TI55xzhdXRWpTHykEp3GQMYCppYA7vcnxt/vpKDHIPILzddQT14gagat1N2VrvB
tT+jsKK30dJkdSzBPDjAJ8UvxbMr61dTVadx3TWWl91KwW2ivqiYO7N3P5ia3rRi
NeIQBvtN66lyiAN9MmPCWP9nl8QBLM6QR7uHXkkUISwOzeK+x8jkDxv1LmCHCsuw
NQ6o6+xWouI3cHrCGuZN/fRwEaStEHa2mQNWJB29/ZYoSOUKJdaIWXAG5YwNuX+2
27V4W+CDV7zOo8x3GIetOmfaw3LS8Hl3KT6tkjYpcKfWNz5AZ04evbjS+BTPYATf
OQ89h5Yxoti+EdDkTjUaepmbC9EhzvUoQRufBIiHOATStMQ47Y0ehYoYRm0m9C3o
xB0uY6TwI+h2EP71T0qfNYdidO/ARro2MY2A6AoFSKRiqrR6bqLYFCn+oJ9Ltlhc
429P4AkHrcK+0c8mleolyeNFgVOph7BCG4oIXtDUOXqEm4yVOeaoXMwOJOLDIKFp
mSPYFtAmPKk90h9JWiJCzu5t0D3NNk3A3xQm6yRhMjoJWwe+uQ+VNsu7a5j90UJq
sDQZER1BtLhYt6+uoN1s22bgA+JhsdOgb/NG+WRmxHvm+yVYY+XfPcFL/HzsyR12
zb0flrIHU2tsxyTzz9eM4XQnoRGHvpQMuzfYVaWj4Ha3lx3F2lRSPd+WAwsi7t7m
Seuozg6duGm6yw0ZkQc2eeyyANiewAcdi1rsMmthMTlm2gD1QK5AuIT5Jn9RHB1D
ooxF77rfRiD1732jwtGc9mCJFVj2hTt4+nTd1F5H/LveoeDhiG2nIbnryqYi4NuP
KtMp5q4jFuPAJd1hg4IxNBcaha60tCPQ3SC/xu4N7+9nB7nKLYlAtOHLAwo5r+he
wAMqmlk4U6e4LocftM+PvqXDx9v9vS4Ae3ajzoWl/5sCUZPer6OvvRqy7CtxYoTz
Ez9EN60hbjsMAXMuDmo9Z82nIbaxZTJStXH6Z1to+G/XzufWTcpqU2Q5Bgk1NFj2
whQoLp1+W8JUEx20EuEIAFCAVOSSgdKRQC2bG1qjBxHRtaAwdPljh3h+0uxHNCpd
RiD4hc2dszQuA+uBh4c9yLX4zs7JkFfY/l3Vg522Z/DBkXX7Qy+/id9xF2S21xDP
AaWWE+6rDoqDOrRMX3F8DXFg1cjJUZkaNHFPHSa/bXcxPOIIp5c7h5Qfb54rcaUE
Es93ZKLvFVMkxDCUX9MmJQ+hYwNxuIk9S2qyAKnUqncD+SmxUrBLps+W6/3yFgl7
R9R7HkQPuY0XhaHlFBcdVDZ+yOxJURwOeewf3b5/9JoixfqPZ57r5IlmPXR/aH7/
Qy4mEDY7OAiFIbjFU7zxXJlGtDNPIrbruoT+kqLqA/p4ocLovB2Za7QUwuj7yHO9
tKQJI+24w9MUjuLTwQtmd3aU398YkOZasiFNQ0VTnaSfjKhBKJatJC+z04uIrMLu
a4VEi5bS/pAwUzs92Ky2ue267PkeqElHwRdliG0hKcFYmFVdPXbecIRCdHhME1DB
tQCRznXwurcTyqXfLj0QaHaWgLElwnWckpNerBr/QoIFFzRk7JGPfGVnQh99ZE2x
PIun22gkH2SqtPOp4Zavw5lhosdO471BvXelRyRi2/PNs+E7CHhtWk1YWVG9G2B6
lHoYMpu+TaPxMu8A8VAk8znJLhOeWRz+gRZfPZsnWIagGYnJZGB1Phw1raB/V4OW
rkdtDBMI3STMhsoKna4jNSI8cp1EQWngOpn0K9eptL/KRkp1xH2EyfVRzCb9D7/9
bDdoPiMX4VKwVlkR4mvQoZfrjlZoPQcwthQ+CUm4Nns5c/tZEekf3jCgjrc4Ch9l
qInlJ7UA7F6h1xQPUR09GXKBHi6xkjnnKv35uXwnN5f1pMp5wVrXOWP8vV+d0hE7
rQeQyRowLh+PpBZYqp3ZHN8F3XTNnTTMBiwUm4Jyekb9Er4ewIzo8TSTI6pEgcR7
ci4p/aSKmjmQVnu+8nWd/rqgEJCAcFC+yOrdhlsDbm5yob2siLQHbPrhi+mpyPxS
eQ7iY/yrfSiH7QfOErxypfyuO5BqkTvT61FFUmcwnmeyUMOR5cJwDxP7x/es+KXv
7eqx0+RHev4WLZvD4U6ZPiBmWWi9mQOpeo4DSHiV0Rfrb2yDrGXYY1KGMVPLLujL
wR0gPl5K2kqT+rMFdb/d8+00RI2+U1W4oFqpmZsUUce7n/WqUzOgD/JtId7YTT2E
THf9rajpeWFPK3nzACuPXtNd8rXOfnfVM7LEvlCvgOM9jgaAWbsHJEd01grCqHjw
kxOznLZp06qYxrKqp6P2Q7aQCG6OqQ/dI7qTe2D9uCTdQp7xp5hijOoGSgHB4Yu1
4SdZwABev2UHygHXRZFpxXGoRqLixNsSgRlrv9Dhug/MIyMcnaXx34KsPX9Zx6dS
ia15qfAcfMOCnaFgJtejd2MJfwdAYWXGNENshJdhVHjRvHbf9sRKMkJXhSQo2gTc
TgFzDdXDraCaeXSpI82yJe49v0hVMfVdKYzWwCOC6gnFm5mOQfCgxyfBSiAt64EG
ufvkfRJhpW1cN5EzEfeWUc9WVrsrngM3dvFxVIxdZshpNUIqDpd6w/n2BXrMIJSp
OLRKm7qPohqkSli8H0e/ihpFzcM7HfvNPIYiL8T9DRwCBUP5qycLG/gOsq15vCnf
1LsMMKWFL8Axi/qFMQL/43nHutUBso/p8lrcFDJTNZK3TiFX+05qDn1YGDdAUA9f
WTBAEPRjjh6qt++5uBYKMfUCzasEdyh+ld58RSAw/1vgocGoQKoDc6kJhfIxJsZZ
6LPan8NjUZTzYQ7Z2wjUKH5siE9XuLpcNsr5Gx4/LfASLTuWVRSoBG7HVXehXKek
rdaXfnS44+baULrfuTezOIQT7ziZ3OpjCVwPgOydHpf2OGaNAtpcMwILFP9Y3y7B
IaF49bKjlycyaz/oO+oPavMy518ZBHXhbGStAC4zoK1gUbObRGJlyArchQE9L2iv
XyUVbd3ex3bPfKUWMF+xw5NA7XlnnHl9CvK1iCbehQ7WIni0/KTBg1wus8pZWEJu
h9YxxBnIrxO9XFcOE8cTTUivIafeaLJFOE/KPGqAmniFBnzUMsp3Gz2JxZlrmPuU
3XGJ0xL8KH4fROfrXdNUOoRZonUK0Ld8PQtn/v/ED9Sd+4GlJcCbGXyQAnZgncMv
EJrLrPgS3GMXKCCRUems++FGk09SIq1iVgJPtEKLf4Qhf14LV3iR7MAQLri9p4j6
tAbHLE3bcloVioNkEynKJcKy+L/2QTDW64ACdo7Ge0fkMHHf5iBOsnVO3F9ymeVH
OWZSnIGJZY+7URCVob7Z+dBNr1Epwca9qxXQ5G1Ocn1Hewdo13AEZdAXs3XdwJ/n
sG0vnE9AR7sLEUMu26cibFqziE5ypHRr+nNNl3irhSm9SgH2HaYoto+fG/5Mppu4
vOPIi+rjEUh5VX06Ebu3XyEFC6rm4Hs9pUlchuvFNUaWS1KdGTZpMZ72jc+d+0fl
XwiAWVNWpQUp5LafdkTxrNFOxtdxXESD5UCeT+4jN1A2mmkTcVhkMR0fHMnLlA2S
M50vDT2//1FQOpIT+Pz/0cZsb+AKesR/yDF9o7zJauK8VGdL5ZFObc5/aL6MIbrK
a+Wofs4abFoTEjitoMXCfNejq/6fN9FuqvnmqweSAVrXUnhLgO0YbPMKz5nMVdI4
angmMRse0O2OLa8tsrVbfd0RoOYIQqspTNcjo/L94AY601MSmPIOG9PVciKTZIZt
bINvptk3RbRvPRr7zMRFJHpWunnAuX90THeHGZa5jN1H2fgbb4rbxa5nyRIgQX9d
n0+RjBokagnrWDvzM7Hc3xblcouJB1U/MkXJQld2R/TG44+pzhS44e2VrXihrBpZ
xAxqT1hfb9vT8WI5rDj9IuxnjY1AOiGlk6t902G4bp5prAK1mv1v7yuQMyCP+ge7
fUx22QA7fF/Xe/dHW9uKhv3ftzXYDxBy+1IipQgn/FWZd5MoNbhh3FHSmJJ3VCa7
fB+e6yHShgH/LitvsLKA5mx/qwgvaLnY37UMGw6w6x76646zSgM3Xff7HEOcDv8d
087SO24g5aCGunIObqjjkPS/Fh3pIZKafQpjw9ZZ7cx56OLQQI7wNRls5L0mTxPs
9qT7YcEOfxDVtfZ+KgNugBXKUQJGsaYS/LMsBJTpv/juQ09j/gjPV9zyRcQ8Th7c
8xatQt7Rt3KlT6yYGQ01b6JMf0we4VUMPz2f02N+Pi5YPbAay4ZRRCs9m69gW8D+
QjxTEv4FIkVs7QsvZW8rD1S7rFCRN8OdFy/dAUHBJkFBDsb4I0oTfgaYvkItYNpT
FP7m+aAnH6uNsPEev7JyH8uymRR/5qW9xvNeMB71jcOqSXfxzPfsW02gXkbAc7Lh
9GYXbGzk8fwyfe+UgB0qZDWpq9KdeOmNMzVjr7kXBLTYw3GujVmKJ6j28sF7yavW
5tx8+HPUpldNobtFXDC1uDkvt3oEuttii4RTgRZoWpUfsI9sVS7N6Tdec5ZLD4cz
jLWBajNBIQDSYImpUxZ5UeUjAtq1xDJ4zugWusAQcRQS2Nyzt93DNBNMv7cc86h8
0uW4n8146VUIjAueaS3R7iVomV4b8dhygtJpPNZE7Xb05DERNAqiU/Mko+IsIeen
3czaGxyAwHtINYG6YZCDrAXOk046F6RA2RfgIYpEwg+zmKu+o4C3aBh4ZxwC2MDH
g02lUiUHEeQ1dMvLBeOsq8xNBj0LXfrX661zjvDmyylQZu6rbartga9+uji9UjXv
A96PzS0lpD2C1DIXlFVj6PXSpIl3k1MzxGTvySia6XtmSTEmhk6n9flSTlADpwsd
TLk5wL3wGHERW2guH2PNkw7V5mvVmLvvaqnMpYlZCCZ8xtUbarcJux3Q1zCw934W
60DXCmsC89K/2qLSHs9Xp4iV4IOnBSb52CUXyTWxONd8y1Dg3k/ZnGIsDvNKjj5k
TpqSicIHqcstjlc1PJlzQVi2A+aYJ/p239RRENJmLl5Sm0fR4cx9URBo6HbksKTX
MlIci+Ho2bs8R9enoupE5gxJy+Mk0O8KEzpx6dS7U7Cxdcs9XSDrjbGCpYxrPEzQ
GfkDKnFTjB+r26vOG9vc9VVi6wGtY3fXfuzIaOt1MLcz4yra8Iid7YebfDqRiPrN
kO6KWgT/g4nl2ZxTWAZ2LDHlE+piUSNbarIwAERrsfhMUYtAMS/Be+XaMGhNzFUg
93z7MXwzKgcS6qKAoCf9grfWTHTV0aLhdDEkrPLnQXjfgJ3IskTACjbUYVyaFiHY
N15M/KGqpufgYhy37GsTvvfwWgI7XDD5UCEbKw5VcHZfDU9MNmt+147Jj6IK792z
nXoV19UeHWtzHgkTkDBofEZsrDYUVZzrEjhSQN/5GjGA/M5imwIOzsw+CiEmxgXe
9O2uB3M8GYNUmAmd666WcRnpXWGrJn9QH/Ew3b6hAIz3ggqk97ma3aqxkWpUffe/
wNBkSpvB8gu38n6ghAHOGrS7Js6YyngH0aTLdzGvCVIf31DjZyii/6MWTdRUucdP
QQT+jeev9tQ8jyCg6Cw36D91BaYkdYNed3hivhaAbJ3UsHbnIL4JBfY4QEKipnpB
T6tdjGZDxSwx9RxzbFG51LieModza0QZW7R/Xv2zaV5prAQ6wr9MlqoxG/O6hvfj
ZfA2TqPRQZrksFuWB3BlDQaeTxY4AR10e9MGBctXqCo8XFa40KS/TlikMUqog3qa
BWoU9XmIb6TLXidhq9/JlLceYgA9jl+wChj1TqFhMYc9LbtU6Z+z/PWjmOHplTZm
+kZ4B8oqqxdd0wdd7/rn6WIQ+t0mbavoS64actXbDwo+PrtI3MZc1hHs3x5QyIbu
pLxlAUTdlV2y/BtXAsmft+/8sTiaAP/au56x2DLrDGcaLRmYaWHAHzyxF4ULmvtP
KMSFCI4Rtwqa3W0L9+xwudQ3s2NsIE0hBnKF+vEljE0hUx+weQE/+rPZZhI7E39D
CumCyQl+EEbhGWoEeJyuJ3WvLR1tCLJFZd64qhKLa8STttCO+2PO3HzDwZTOeyzL
NbUfBZRY//jRZifnplRS+Rvp/d2mrHXL3S0VEK8K1auWxSbpxzaE5dlbgfRrODDo
86CWPfkqV4Q2CbSsbzm3MNKiSgFu+l7jTDE0PJk3RMs/B20JI79CFneWOinQ7RLa
haM+pla3FwvHPHR/FYNjhyE1H1aPxJVh6oBKrsvIt0eymagd01+JE1lNtGatm+QW
ouAf/dHFqNCvg9r+mUYJIet9EN6xUewnFzDSOc1n1igkBlCWhaquFjNS30V1D9Hw
zr4kaVlnaA/TotJ09Mgz1YSbVUzxC/4J4lkeeXT+0qn8s0mxqoylxMV4wNxOOKVw
KeBkhzHX+J6uRR5O3jQ1chjXuxtnwtuGO8PzPAEpr6s1SbGVdFxNdYNET0ZangQf
tw6dnk/8+27XrijDn05Oy84I+ovSxOAsX6bzAxABs7HgjanyHSVSyorKjLLLfpVf
5KtNJLDgOwmeYsNs1mK+tbTx38jNNXpRS8TS56xtZqV1TsQUxJwKVZOXhxv5xwBh
fcwKMrK1Tk2pGBF2TQm0ZXRtdXnZ5be76h67Lp+bCzaasIeOSbJtHJ9hUpFwe3Ee
Z9h2V1vrZZL4nIIbxb4hxXpc4FWQhpkuLjzXr28SxgnVN9qbcL2+ZzfqrsftgEQA
gpg64RW7fZFTvhRSmlhpiTJDoFYffLQV4xe29a1mGPoNUoTdwbYC2nM0y4HCUNt1
WKLs5leK9B/1zcCmy5ZqypL6mLQz2LhcH0ElzoZ8oEwz0u9NzSyXNRGEFeGgPu0i
u8CfZtqcTk81NOaGhr6UYkdEMwuL8iLAtvYuqq8kI9Mhn+tbOjpbw4g+E1OWd0N2
LQPQaDJlJPHNT1l96XVJxTRLr/fs8gViXUxCuNYxFW60cPbJAd6KeJyZgCi+rhDw
Un7BBvt/WSDPhohjEsEdw9qMerUzAgyAApfebNiKkq+UdC2VT6SuNyhNLjZUFdCk
b0RJ+9C5yv6zB9EzpAafMWyTi4poTLxKkE6kWYxZF2TQ4pCYfJKyN2LJkjeeE1Gm
NMpQSqWOkLhHDFYj1i7A8aeo+0tIVUfokNuFl2Cydoe8KRrmFH6QF8RKKz2eemsR
lyHZuaRgHyRSgfpXKRABTULcLzd4rh4QG+kgAXHxv3OhExgUE5PvT893aoAXPBQw
vC95PCdJ4RvIofdt3UzLbXIxvtKVLY0xSovlSpBllYI/qIzdy95lHXOxUaWjRhPG
pWABHX2p4QvGOadaQGc5XsI6hCvTmpSg//utz2rtoCJzIpeEYFKdduGBdJplq+bK
hBuHVExZlx4hCV9stTueflh6re0eiGahOnJYJtdAGnDH0wI7I1+XZ8l2WXhnUq4c
SEYrSdRIj9ogJjBGBpTb/aw/JFq727fq9ddU3N8mhyK9lh2Gsz7g6kyr000MZ+H6
vGDZN7NyPt9SDI1r600VLXR73Vw+LAEeS7xU5cXOOBNUIRYsvTUmU4nWFT6qpJjS
bb7rDhGg3jbBN9YEh0G9NNPd4rmlFfiM/MTKKwYnYpOpUSx7i9Z/TB6fOcdPQ2Ez
43IRM2TszuT5WYDMmzMDe7bglTT2mx+PKC/PcU596Dv0awz2mXTdFXTaNii17LBn
Uwzz8oSq6YEruX+XDjHZFw7o263WS/3aK/25XScKRXwY/S5jLHNiU7coIw7ZhuaM
eaiNAuk9JPNjuofNAhSRZmlb/KFn0wGZNbbrk3vJKN+EZeKF2qNsAvyzo2O6me9k
RfClwU4avN+ko4T7Q6caHqkA3nj3ujpZSY8/m9kTxGu96ja3ljOFIRHTj585eyEz
q+ymX4DPajaSXhqitwM0gF3/XSHaOWbx8+9Ciq9M2J/ZI37Qy0hYliZTWMFQ9ENl
5uU37wQrtq++EHRVSHYqy/rWZKWu3JuZWTPgGhNJcCy/9Qu8JJobd1YzazsK/bH2
upfQxcTqsNAGFQOtIIj7L61YyAa/LCUUKCVvklRCGPvyx+WcWOdoWuw1saaektVU
8d2ptRvNryFngAcuqm4DpW/G5VNxSIENCkUOw93ToqWIEELDBkBJAAP1AuhJFUle
ABBbNnuwt6m62T5g3q2FCYBM5ntVyK3HN6kv1yrmtuhD84MvTgBDBIOD28SdwqPn
gaRREW9ERV1xCqLuHYVTgJiFUMwwNeyo3VZop1aNzEyqyV+SMeGao95NdT2WMzy5
xM+aQkskDHdvxGTe3M/yz0pNC/KOpQwGjmeO9a3GSL0OqEicdbsKlAqxQW1dsqYo
jh3aeodvroTxzahBVpRuwBnPCBXz81ZsxIHB3b65P7dQcLZgRxikKdfsvWnu+HlX
g8pZGxkekZfMQEepLVvxR5zCF2sIAuIgNVEn9jux4GEikRxGgnwoBk3S+3FwyS6j
mLamR07jD+JtJ0FeoNoy4g0yxejmi0iIA8dwLMtUozPQ2NOSG9cIDSF0MRFOOGD+
RrtkQ579SGaG9SPGKJ0T6o9rcOsnOOsUb9wZK73zrf7UAfqYK1xPMdWJTLRM6ovN
HlTl+iA7Hgl0rT2XlI2Nv0nMW/del8RZlXigpbbNNzMrH2OU4oYN+NppFDjg5sJn
6yKUARJvk1YTwm+XH+UFFeXtGA+YVPlNC4K2g6+MbID5u7PVomG0IMIF44NUE9a9
rGmsq9IHL8xnpxDI8Q9uwEnjpwbr/CPbEEcPwPycOh6+9vLHzTV/Sl9STIF8gQGx
SWq9ZKWmMoRciQJsQBK/UFn8vr9oyTU3DXWuql/8tAXiYbjmP6vy1NCwVWbHAypG
T6VaXFMSVxjG11Oks9bpHZ4rv+lRHDyCLa6buoMWcRMaO1NbjHYLS13VYVCX3lVa
A6tAYUTB36a2mhMnKMqR2rPlq8jRLHdKv2VcymGNJ9zwcth9oOxTgk9FjHVOo8+7
APOUFn+BRzejK3NWv48StcIrQQ6Yxm1QXzHGZpZnqLnqFkqrlpigc08oRV4m83sL
CN4OPGJt3gIXBAWtSSGfM13yCLvaV4aS/qXyCZkhdUEp0vc91QDGTkuN87yIOpbr
g7hLeN7S7dLvYbdw/r9OJjJQpsfVXEdfJbzxIvyRlQekR/sG0kXT5/tijq+uwvAA
nXxn72CsEkpGppd8F/gV/GrPHbCtN1RJG2RwxZPJM7eDXgGmzx1dweLZb0MnG4uL
IolDu6kQQRqgJdzFL6gq8W8J5GIITOMuwuE3KK0g2HqoFsOyrhHrrga8gRV9X0DV
Uy7e1bafl9X8twgJehBL3VQKlXXUPTvMNXWRjhLSWX885R/N58jqLajNQbMBz+EN
9ZFpCBEDz0kkIW5euZj0LUsHNAKqh564eNwPG2poz6aUVbMu2fCLOLhJmA4Qx/Po
z+sUB2TWl6r2biZV5muJTxxcwZ43mUFkw+3+tsZrPWpfV9I+/VXCEVwxuoDZBNno
Rj8EeYZu3Y8t6ZjdXW03s+uGZ19WIR8ExDZtIdgHLflADRtSsaiyU1IzCo69NniG
Nqb77lPLGatW4Ox+JTx3J/Z4AV357OdmwdfJ1vNXbWfqxEjrkjcmq4+HwI7fCBGj
OfYsy7sDMMY1CMU1Q0L+NV68UgvRovi2Oj+6Ymj5yzB82eaBBVGIFCSKrbgH/POi
FKxr7LCB0JmlKT0+LZIVAyuCaVTXdvzbPbXWUuG4W5ZMV5JBbKwfdLB6eO2o3jdL
R+99c2yipB1a9ADQLmdvEa+HDni96Wgf8or7OqRzq+NPs2mSrYM6ty2rXtouFZTk
OGZt0wYZkzicdfpY8NTTIs9ZeFQKoA2X0OtBT1oJkU/UfhyKwOj1z9sHc/1rAB+B
OP81IKC0S0VKYmc7bcTqIpbheuMek2nLHEM3twx53Lww9ojPunog9FbvaB5lIJPT
DqRFLYTWVVs9LFTWhq400qRkkeRO6ONDCFnmvpXZW+4DuBwAJPb89xB7LQwOArpC
x27oTGH76q4WQly389xfzuGtfkR5MXR6Sb+hS30iHdj3f/P0SNiNddHAXG23VAUZ
EOxTgZf7O/nYQDjbyRv03LGpDpSVy9t+4NMZP9ARyg5uC4qHUSeNHnXoK1OdSRiq
Nacdq7Td5iv94b2zXpiShCCCTbpm2X1PKk+iP7zrmLGQMAGovd8ZCL0LM9mKGfDL
2ONp8k1J811+7NxYcKR+T5ZjfeaweVPJHyv3JNw5kx8SiKcptayUAYCxK/m8d8oN
qwwbCbAn76j1eIubGA2ytlpiAnY0YlN+3m4gQ4sCQ0Cs4KCWgCUEWq4xh+bI7CTa
LJGbZIF8Urk7YOmAOiBXCavMD77LXL87T9OTsR4jFURYrWUWqPZi5LY+h+FVQO8V
/dSaVCEEjlGdWY1iha1Gz8fzZTMWlFkfj81bf2WVwHAET+jErnZF2y5+tKaQZ+eA
ssO3zozgaXWgRBv9u9Ze6uaIBDykbbLE06Vzjp8Aj65tp2F0KdR6itAo8Bwj1rgx
da3ixeCWV8nqyI1WSw+S5kZYKs7dyexRecaCfMVZ62CSx5/ECNEUGNigCFknX+eM
ZatsYMxh/dMalFkg9cqd6/fyLRshrEjWqnbLhmTU6BuC9QoBSAo5hXX4fsQXdy0D
JMHMxB2PvGLgIFcpppmLdukDkU5Xd6geoh02MHgO65fqhZOBvisMFRwahfUn5mpX
v6N965LXBcBt8h50BOPNDCVaE/Uo596r1J1FpgmJPoUIrZT+08TLQNa+bisIFyIJ
3HnWJ+WXIJylzCfbAul09W+tcLaCMma/okc02HtSSnKzSWzmkfTmNhAhjr6UnVXn
tu06Exj7DTO3AvYlAKJ+4b4KS/Cw/GIVwMDb4uPvVSZS7uCr1i5WtRimL2qgyorb
IUa3eJ8kQ3ENb8o75kszz6bZ0PnlVqKQnKPMfO8rAGISRkBsMnZbNnl1/Tm2P6tq
GqhbKSney9plg5X4D4z/qJ+WfI9GG/wME+Lgr++neQo1sUqK3puskYxEvgNTuPet
jTVg/fwSSy5HZNgudN4Sdi5bPR90xLfsef2VVn8KDsxZvWA8KYa6J11ptdnFGhLI
nDMnUOZWovrz+3LlTKgN7wtQPzyZvjt/FxwEb8swPgeubgQWUZchjDfr5pulUddL
Vpfr7JOihZMTWbMWnD4KX/+N8FOgqLfa2yqOsQgUPrP+nWX4htexT40eWSqQpU7L
CHAceqTfhivjXOjz5tPV8J0Bso4Lg0WN7LYNuI+Rb17/HxVTCM2gFLjBM1RRhRor
LrMQgUHmbfqDCS4gmrkPrIhE4vaI6FDSbPfNDtzX9HQl0DoT1RNvpCZQWQhdZSvQ
Q6ecfGTSzFnKEBkwMmtPlQK9LqHQ9umvVy90ud3IeXxKoYfi/BYqpCWMZtRSyZPb
twIG9IhUetK+zrQGpASwsd8F+kEviKNkDhsnOsRS8vUgT4hmguSm1kvoSFf18C5y
qrgNTan3M7EoRw2LVVg5FsibmrpshwYFm6P8zicneNqyDO+aESKbXylTBOMl8zMu
baMn3GBjFu8o7Bp265KzzmtmQ1vuzeVEbAsVtl5pbR5/73QT0N3qiVD0z8Qx9K2L
nW5edS3WQky0a/b98p1KtSLLKUlVvC27rapwI3UtREqHbhDD8Qnbe+CMtKflT+ay
3JszAajAJvLqtucIQLX7Aa0Pfdogn3I51ka9tcqioiTAAi+OZZjxIREBnVPr6JqG
e1XvP8h4bPFQZjJFPqqvOzSQWCsbzDhNFU31QJYXnaJmVu/o5zM9Wv2a/p7AJk41
IDvAKzS4qJ/dF3Pt8Ugn07Snn0jywu471xIYJmNIy7oGBpbRJUTWtf2jgaRskurr
Kbg7irhtDsGuPP8hjNNCVp+69YRLb47mRvFjotSaIOKrw5Q8MLYqSlCuaDYpPNTT
apjs71/fCOhye2I5zkf9pJiywQE1TU25L1A8/Lt3AvdGY38aVgzWedgBKfOyxwJ6
+SNQ8OF2Sk4NCSoQg33BiRI2XHfIq4mHOlt9XoId2KIhvIfuKwTOkQddybPCuohs
Z3szPEMQF3XL25KAY2aOLJbSokLeZMtNww9zpyWHPYjvCb/2yYJUCPrdGa/Gdn2B
fNzKMr1O9AtgoxL/6FNfMa+RgNvY3XesBSnbVbey890BxncZ0LYeBNzDckzo7+78
bBCl0nGtD49F1ejuc5dBITMSGRK4y29AsCd6KSc+PV76Acb0i/35Mptdxf2/VGd8
p6bti+JIaUeSaL0ZGsvKMcSLdlqGr19yigQlspDjbnRI/0nVf3dJwJSKoPRq6Gg4
dnFn9HzpdMoDgw6AlZ4Enx9AfYs41xwXBga9liKOd2+FcThwk/SGsFgBLszPmuyb
HG8jMsmE+2qhe6zPP+bqa/NY4ouI2/TRRHhuAQCsRBzAP8UnLkUn7TtSGXwpQlHf
K1BLPOVcfoq8/lWJ8fQc7tSeYenbpAhovYfXy3muI/yMmuIRZDYOt57ZYbavYMWV
eSPBC5PpdY7LMoQVdMpx/ARiGr9maFTMtR+o2nHZreiDE+f5o32JS5YVRAh2Gxj8
8VuNaQ/wA8hLNjyVh/7DB0PeAuDNa96PScVlja+4ks7wbGL28bbuyWM2ocZbzGmX
3yxt/ntYw5F7ElczY74N3a4iNZsLO6G+DTwHYtMDXrRMlT/nDng51wsSiFertWh1
zWOEE9HSmgWGuGcs9pow8Gu0TPwXSnM2iMrKPMt/EOJEl/t9kL0UsAZSzaRa47iY
K33l7B6J7BicOSoOG48XPpwIpKlFje6pKUp8qSmjIjT1cZ/9ytzydLs4eq8Dng7u
/xyxm9KlCM/cPGrgII1WcQvo30xNPW2vXk2q5QBkAKYR7qcpwshaR7ks+vUWccT7
a29KDDkVSS75RLTdQ3TLopm/e9BfJgG/SmsInmjL/pmn6gtuAXPzmcpLbKgVvVsM
09Azto7wQ2wI0ne0Z6xUAFHJURWxffNaDcqcKse2KKJQq7DWu6AswUjIb0z30Mh2
EpWAKGW8EksKGDw+KHUFJyh45oGEYR7XM9ub1fwviW8l861W/yFi7UgHeVv/+zZW
sf4LBG9+MBYEyjHfwyhGQB3ABy35KCqy//pZ+aIWnPReaTpux4+bbe31c1Q2Pkcl
Qv3xEsWip71ipnYogM271aXrDFBejrKOcrZ3SEgDHR6PKMyUG4Zbfnr4Wo2aTwj2
7MvpzqdvJ64A3XFZjaxBwJqmB8b6bkxOJo2cuaMLpzHu19bBfuh6n4pvOjtjx8Ac
y7ZxjhXobXWjRX0yfoFaYCctwTWxfc+7Cz42z0cyUqDHN0H4VwOTtYLPUoyMxkzI
3GUsRVuhdsJ3Aawi46T106tdAPlF/RTsikYvgn8oU12arTsi/4d5deSNaoohEGqB
x6h1HHTvUjCWUWTBPc9OQ0dYFIqSldKmO+hXewGdcwgfdC3azxO4Xu4o0Kd9juef
58rIb5GZkJUEipQp+KhUs9MJbz+uxQSXhjgmvI+ZfL9KoNuJBsByDF5YDDI38Ucg
HdDxOLbgsrfCf+wqNjuSFF285258hmy5Dv2E/ypYZMTwS8B47GjqKNXYa4Nv7yZg
yC4eZk5xEQdNTBYPlKreJ7JGhC39KeJfgegtnV1eSGdETD88/OCBKAzusdooiNHo
Ojuu9v9tqyVb6X7gKCjOdHO77rhfb3XdTfIhxT6OYOP4f90Y+zI5lvlSK48RuV58
owFtWRS/ZvQ/sF7RlxopI9JQe24stHu/YdgMDmDUvimpnftENZmNS8r6MiyRPG0i
YpqWJvRvfEh8qMY+sw2NGfq3npWnQucuBtIkgWjK0+j69on4Zem+SnK/Kl/KHedU
qGF5FcvNcKumN/NDVcb+2AL7B2iaNbz6mRN6m0mNGZlopgEU6nrjCDnmor5NhgaJ
smSd/T4rAeP2O62HKtjCkCILEKdLGD0ztT0/fWsNw3CvY1nh2bWvl76a4TnYp2om
lsk0xS15ml34f/VoaV8XZs/I4WZP4fPe1RYrw7YPmnbIAisA33Fmr5q+sOZuazkN
9HGVP59NzDMshjHade8uhT7gx0Srjbs2yEstQcPzrZXI7gOt0s75XXBa7bW0eePa
+/SkCyp80UbcHJiVUVJJ0Kidif8eyB60PYDL5lPmEf5YLfVJ9Vrvcbm8jFeAwCzL
xfNgIfXl/EYhJYixgb7LZNzIBAxnpS655dbaC2rJ7l6IGpExFbweohnKRSaixSWU
i95TzAC5dLLiRGjSSWrJikye+RIN544RZhLcFpVe2EwAEV0dCbmiwzR2SLxE+K2q
EaU7GVRXWb7DeI8YhNG7jL8U9GRjbhr1IcccgcB7XjwvJ9mtjgIU6IX5WN1IAi/X
ax+AtrIvA9Xi1nmcQ8U0QgGslDEGKX8SIlhW52u9I5gSrAKELYT2YiMQwEHiymIJ
J5UX0fsVMgyV/WBCpde0DQV/7J3IJ7HuS+RlDUfVPnoW2bMvaZDIXnNFD49Zt0WR
qNJBwm3xoKocTwckWDfXAqdNv0idvzujb9rNyAEBAv3zCUflvCT2bCOdiuIpg03v
O6ilms+K0PwKAlaxuyftlyy6As+YpGHv2sbeislhYb7aJXNBoYYQ6nT5Piamp1u8
UvxAiCSlLRJhi5nMXnd3F3wRAINHDLMzyN5LxQ6Dd/MaTxBM03MhHhjz/dtgqnr/
Y/hSwqEq7r+Ly/a0xCtT0E/hhCIq2x7NDjeT4wNGTMb4fVe7teu93BwMPJiVFFo6
sLsyHEYsw3bIHg6a5vXlk0XdL3f4uWVWIG9JJPjp8m6zkgdFYHmMDkJzj87FYD1u
3AriLnSI1XZORi+wXif/bUvlxcdRLEEN7bPQs8DoxmMoTonrSHUB5YglqaYGVqA6
YLx6qEf8W4XxCGwGRn5Iavf5BHstTLhj6zFDMdl6CTub6bMP3ecSsAsN0b1IUZ+w
DtXL9XHU8JKowBkpoc8Nm2Xo199pj20WiXVbXqKiYMJb7cCK4f9LndMtsMAh4E5W
Oro9lPC1S4TnXOmOkEf9ubpcLU7VNNUcdclqpOO6QFlwZeSkybI/Uj8D9KRRU9Zs
gRbYiw34wiifJo9QpIq9GHEXxhroF7qgPR087ldzlrQjV0iABtL1jtrmqvymR7LM
v4Gdj/9PWewM0cwyNm0QlK/Jzh9HlYGuOdLiyRlLh86dc+O1s6YQKfWKco3Y/vgn
w5AZ8zie+fXhBBK29T1Goep8eTPy9oUD4pYfw9njjeTczgygLv70PjAVY/VrBmLu
FHFVcPtIIZ81AL5sgwMbB1h77uB62fa1nUTmu2t1RrD7ai7vgmxVTim/3JEp4v4o
f3rf14TdtLjVRFoZyyGGofPC4sjER9qxBrDfOuAftBtRtgs+n+hqyY1zRVEIKg9u
2RPCwmxyXM/cRx4v3L5yszIoRaoFE1PxhTygwNiV80l/DWP4Q0I4dFGC0qQoAMAt
zWCy0MjoAW/y3M9/6Bg7ry+fgAcgjiBryvQBeEcewZjBgPGpgzv9QfaOZM7UsijL
bnEuWWPuw24Kk5lpeiTwBgaAMoyjWqihU1lFed1dV+YAxM99VpBo+OswGynJdFJw
zhFbZjrAKMYsJMLZEJHk/LuWf+UHhhXl5UgjX6ejW0ME69rrIa92cLc7+YRAhiJG
k83C30suOJ/1aZjLKtmytihQ6HjD6UmdFted41k0c/TQxxz5l2k2cB21v3HGVC5h
CxSlBfd5MNQ08Q6cwGti3ZPVVb6X6QqSXegqd+xacvFYc3AdBBLpP750c4CcVxsU
Fy4UDGPgHl6Tk39JBrrQr9DsLOuEDqJPd7WDR2LApdK/864S73NaMXY2ATRyHVXG
y5HrcW5Sk3GEY8YQ2DGzMQkWwWv3T5p0Y64scxAiUAofziRs3if+p/ZDCz4zj4oY
HegStTZvvqtgokiF3XYB0IXaFDyCFOQUh5cyKHpSM7LnsmB+Glp2cpMyUYAGRmqe
RcbrxqvjQny8n39d3aDUh0S9j2+b+02NKLumZZgPwVtCMyJgcLs87pY4SGyezcyy
lIfRLlYAjqpomZX5B/iOHYMCt4gkNp0bHpXtae80glBSlOuBQXnN5KiQRkiGwiUp
mlFg4EgaxYHs2wxE72xBw5weeORZjWXznECScMCZ4atHB+t82RgJaGZ/xii5SUJy
tJsCqlVCgvfXNFXp5pH9iwdnBkb4Rbp6FjVvSpll5RI4dFzE8D7Cj30KN/btDDG+
9XW0VjxbWgRFtqr7iiLSETxku4URYJ2YwxGR86BpA1OxpCNRNCKJMIZs/7/flHbD
ZQNdWR5FJMAGyIfNtp1u9wN6Er4Ynp7ZHzXrsz33AlF5b0nxpsZ6H28ZFHDHFhlD
QhHNMcvZAHgpVvVKAaOxxq376+JDy8/a4LzFNj/CThLx3CG/R/oExHxytf16xTL6
fkPWPtI2WW9H1YRLQRYlL94RvWDtUKXsYsXc2TDN15jSJC+P4zHXITTlQK2anU+W
a14z61DCnrZyma2i4KFd5gUnWdvOPXWXLx4h6MkjlM652E/sf2Mwf+dO/hDYFHjI
DD75hq9zMrlnzz4F2+E0tg516DoEVHCjGji+Ck1GhFwxdQLvt4Z5YPLVrq1akAue
82iHQ0xfvwXKwCxd3zeUcnqmaHJVKfV3+KgYUcT3DJCgJXe2eUajyk8edsP3tWF3
Zsu/+FpEvvAQ5U0H9o34bu9euZjR9vGj28kKkQ5xTdwzP4x/rT9dzcnhC5I3DEUC
Mf8H5wZtuEsNCAOt7kyTkd9/sjKekgzB+T7QKO7fUEsS4XIzHOYd0GfiZr33xlrC
zAnoYnndc92wv7yJPvVAnXyMY8turOlRsgxgujbTRDktQj1qELZGQSb7ajFIcuIY
1u9TpK5w7vkFpuYCVEeLj5briXhFqIfTRhn2lS11WdfeNCAZ2ban3VCjDxl74zOA
nnzV8OpC17mqAgQqW8RectpzyI6Uvw3GPMCKC4cHUBrKlNgoA4K9bI6SkNgvvZXn
8UiBhTuuZTZjn9u8oaUpoWXCPg48tnFwaAzSxSeZusUVR25xZIqY1I79HZqa/1xr
Srhgmm+gHm4I8BylKEFeyVJZfKFD1eFAPZ25s6TLuHlfqRfIvS4Xo5cVRrBojTeB
Oem7NotDfg2okv8objwd/CNIS5Y2RYRCP0XW+32Thm/sQ4+6DD99Y/cD8hSwH1dO
lb5CpLHEINIbbdzjm1W7kH9ewR5g+D2aCMc5wbIAKhlyPPtQk4u5s7wkrBXr1tXy
EbmldO4DfqS/GM4Y/FJodeTBg2bMvWm3fGp7hCrjysQClJ8XEXEBtrDbonl5h48r
82kaJkuNwNQBmogEUl477nZjaDyK9y+DOue4VxUrebTOIad540oWwIwjZZSv6As3
pyapW8zAl46EbvAXw6ZA4bMR1DBoxSQE9fL5zCgmDBFqKK93rj7LvQ+SbNjeKGdT
BfYp+lHZjMr8ZvQY9gXuKEcqM5+doLrz6QpBkV/F4D7K1ZAASEzd26uAAM6/pMSH
lLFK8bKvI0kG74hBl+5IrQMfwBbcXh3Plj1Fa4xBVGVcP76FCtfEnGzsRb92qntG
9YxdaMI3FlUx58I1E//FiIeOtdMJMm+1PDO+B7puCtmayPeLlh+szCWcxlnmYQYg
Gaf49yLyEbxHOz/rwMtD8gwMMOOT02lHf7rx5TtvWSb7F1gX2XuCqAkiyJxSIDi/
JiVJgRVNhTmIEyNqkqxk0o/D8i0mlD5DOxkGZnNxSPUEKY/ltyKRM6v71xt/g8h8
oRgXdd4DJ89X5eeqKyKQGt4VugtwDC76ybWll7k+wCYxAWsd4WQqzghWAlqKU1ka
OMaPJPZplcD3xShEaZNwxIOZ60tqWHLjo5Wkjmin2LIw3A8cG/5dTXbKaxKBYfFU
+zH5y2ULfUyT1fuheQ2P1Xcv1ScmxLfp2c03j4/LE6V3TzZXViU9DR5sWFYUvqcv
nnVnAEZgLuqD7XsyU8bNF98NX3llHuLV7cDCMkvSxiwgjpALZoq1MQU8uqxtZ42w
NexBXD+nHZ/ae/LjjgBcFlFvg3ExEy4QnJ4+7aog7OZe1f2KhslQyFlV7IgOTZNg
r9hPAwMf0PFbncSYvsQURswhrnd16nyBy01ZbsDc4iMXio0xa9tuRoGNEQEFi6Y8
pqXb9e2AASTCq6Fcms1cAQ4ILvfB7nEv98XK/m4W0tYyzCla8gtzl77QkB7WC9H/
zx1P+8A9BiyHzK+DFy8F7zp7eyzp1sdq8r8fug0QrUvvCEHDmVN7zatEwHypzfiV
LiJx8OgTqnUUU21LYftsABMYGXFR/KjcMmMyxeS+twAe1AJalX1pYyiOgoJ/Ispq
66uPW/Ql1HZPnMyi+laH3GS8yg/yst3d0zGr69qbAb+6EPSF7uxARTKYWf8k169Y
ANIO03eui5qaV04i6RQYc1KfqJPDUPACdsai60vgDb6uMD6iifjBpbjMPZNb7Rkf
Pqu3zpPcptP85NHvvNkBF973ZM39ODoStuJc7ub7KT3akuas5Q/KPvf8N5K2LSX9
xT1NaR0KDWFxrDSyqAHRKXvYnuWvTQIhljFHlkAElXoYsHATt07vYwArOkzIkdZg
Jk35phdZ7Mnfa+GQEMdNN4yjzQPQRys8iJFNPPD4syZ4mCksseCIrYTrvWDsIOe5
KJy8EshY8VunA2l3DX7y8pndLuunDRcAHljVNpkgvenZBLobFt+v5aEaUhyVlGWm
VkSCqmLQddTVkh5DTFlMDQdvdUTBoMJyNPRVsYHNR2OLhb6HwCoLnTnCZQ92HHyY
Kb64uf0kah+02drfxwxmZxz4ct3TCKH+iu2YnFl9nA2kAowqijR2IO4HBsWgxll+
VDVCOxDelvTM5ppa3qaU3lqwfP2bszFUWUHI1/pR6BpLsfM/7MkxjcJCU5gIj5td
QQZiCIzcJyI6zOrLjJvJ7S7AOoMGIySQLyvTPR0yxt8ZBduqzgtAbed6fegCxpKa
FYhMxcPvGri0jHdYbiACayfI5u02b7eRKEm0z5B1MveFD+eHyT/zkZpQi4hb8/R9
oKOgjSfcb89lveA1KrEj83aPVQrUjlwwnN1bwXJ2OV0rpXJoCHMQHi7nIt+aHicj
ScJCQ/rTFmXjRx9SHQVCAT9uN+s8TwdhKKn5lf6JD5EMQTVCQjlb/1aPJ4/mnYD1
gP0uZpPPmW/szPy7tNsOTm4dd6j/7GNA2raEZ1FYpeazrShxSE8qNbzPnZSUfn8p
mLX2jnC5hfOMsRrH4aeVJsGIMTB68ugKWKrIzBV+j0O4HRSINJLhNogHpRDmOAri
Oi22Tf7JW+qA4+eV5AWE3zf1C9jpNz2kmDexPCj9PRxFLkbCyDOgeX3w5BlnbyCk
qtjZyrzh7YqshemfBvtzCpvSrUnd+6AO+u4fyMyLVYrtakhCNuBNebPCq29iNLPR
kC8EYHdbrjag7DD7NAeyHebDynrnEuzR4Bpj/xkxLGVIAvTI2OHuYeSWeqAdicMw
Gw6fZNo3IAHdcQNcl3EN/MfZOUiLjKHTBRZgwanScZgU7E5mqX4GP3I4kZSZohL5
Us2aPMv6Xt6BTjjv7Oaynor9S7j0j+a6SN60kA7uR0zcAYmyEYrou9FuskMG7Cwd
a1wQMSO9cH4qBNHtV1BF6Vm7kymIBu2H10h57b8EWZEE3VlGJ1C4CHCSJkUsG/Pm
iIHJiX1WvGT2ebVSRBrkn1MCnAgLQTtwpB9sBAP40yq+5Pr++2mt7gjvXuTnYJMH
yjDnUU1Mg2OZk+HmusyNAaSJu7T2vTuIyIm+XFVXpGz3UGLnkpjUNHI+eGg8x35Z
wsaQkDFdV6LRR3xDKz8MCLhPFRb2Xvv7ofWGLj506RoDlokbcILIgTLhM0CmT6N9
3W2xRKwpnMhxCOSvFxFSdHB0AkpX5NQRlDJ55YLehOstI4Sfgeg6p4F9IFXx+ROd
pH///GBsr3Wxf6T3Spc7Rm6fivaRUbL9ulxD/NahyIL+RbYD00oG6148n889dcrQ
+EYu9AdYXqU0GWyAB4+X/Ebo4VF4B+nSC9w4g3g2vBYzU+azWgJuXyWdE0i8ZBgn
8RCws1YWiuLngu5uwCOAISf/xvO/LGqSEQ5t1/sIgKAMM8lF0smH+VI8VWe3eRW7
0elZ5C8U1yOPPJ6NasNaFjSNYtO8NpROLPJ05FKFvIoAnbdq5V02ZxvITqeFKqvk
zdYskDPtW6ljBOpnhkM6kBVGHaRgU+mu1hqPREOEx51Qa1+kcHENP7rGIdppjd85
eaBmf4eRPc7EW2RcLxHDf+OPqLr8klMduivTQMW3r/0khUASIIAu6zihUcmWjo39
n8iaHGGGCOS3HKcFINCQlVqn7kAttVb/9e/APr+5EZeErGDWG/1NSh7TiCqYWDFu
/TQKL+C3gYDyfjtSJoh/dD4BpQDiSw/7LG67rYm07Tz0c7D5ki6EUIFL9D/L7ziw
GXTqeQIEyUSRzcc5UHwlc/vtXXejMG327zqd4kTw2Mey6EpiI/3k/CfK7BJjcyNQ
e2UN+ydEiT2Ypdj8khVBpaeZKm4Ja0TfUOE+sHDIh4WrXrvcbEnrjdfbHN3xjdM5
CnClisbRLUu3LKGsYBioQKeIBiSrjT8COxP8hvdpKPtpr0HISBu0//dWb1IRjLL7
MXhv2wEMmiK/4NWfVM9Apl/K0jivrDFOoLvKAMJ7K9kshdldkcVOJceR2i2fiA4A
oLQwaCm4/IPmFBc1BSroyjMuAeYwgxP0Wv9s4h0BQcp9Fi4ow9dRg4CuyAHj8X6z
nx05dwDA2whkbZ78i2TVCGi/fZaM8oVaG5zrxnXGtHgTOA4vxPHSn+EoeZbDJTje
K3M92hnHeBkfin0sf9HvzjrV4SSzlreN/GblGEWKgH6SAL928kcSeNcf8rP6TEZJ
JCnQgWI02LMmaCdTqrwr/8umNhbM6fEEG+ov0msoXtAIcfGWqg9TyYGFsyjR63FB
FHTBjPaKJIVW0BaiWSPinja4nobW0R+5XAtJXt4iXu8ybA2IiN7oDUGzRCKlQkSP
Kiv/hmORUYvci1cXrKGMU2CMw5COc7w3ZCJrF0BWCRlwo6DiaaEBY8MwvQOxi46L
YJhzDaQCsabmj0MhJTqhcgzjQgx7VhXlfnGPBvqrewqx7u5zSU8C4eh2VPEVUr6q
P6ZwFASuP8xhlKF1Aj30zBMrnohZZnf7G124z4Q06q59U6pk5UpsHPwyIeK7ddFg
PVEn+zCt6YlCd1m0VUFoGEjWIW5eb5PaTAOf/UJomL6Q8sCW9uNQ4+5scwc+4mxS
jyZf9jHH1KmuLFZQlv4PfQms9HuT38BuTN3NdS1Lh58Yv/+rBeAbibIhr8+7Dl0T
FamksB1bcxwjlzfWZ6zQ8xen+n0i25JpEz90e5zUQmTVQk1JatyQ16jaPsGDxhaW
zzolK2t/+Uxp7SBMFS/eVqxNf8KeRH8aYJMSRp1mpWqwFoMVtykbYCGQgVT+4E5c
uZSi971UpmHnyXvrMKMpopVUuQnJr6+lcl5p/Oh1z8cqPEXNpgH1xSE4o63JIimS
s4b3FV5zSFxmv3qBUY3+2kAuDbAT1SycBKXdQngu0W1J6xQ9Q4w94GX1n2kDbFzX
Fh665C0/qfCkXVj89pKonJFh6zEYAgQYaWxB28cTBk1us8yAho+e7R4P9+STOnLd
mzA3ST3wxcpzW7+DET/eipe+10mElmoMT60UnTZjjGCe59UxdTclIIQPv8P5/V6B
bTEg6a1fFWqhQc1aMsdiD4pxZ+Lw/gKZ4CUvHbqCsORUhhkrvBdyIlnbi25R2tLz
c7A97VMMV+Ix/wiqzgt+E84SnGlAgWUVxEhNqMZzVwaeIcimPAEncTnEYXDMLbwe
5NjSHFYSmzcOwZTlc3fTBq9cr9hFt2IOFJD6kf3dX91iK/RaIkkQVlI0sZxZNTGD
inRODHkOGs9hEAea6r2CiOe4mkbqujEkH5z94A5KOLQD1K6lAN4t6fmbPRFh7jjK
mzLeVcNAyEcAzbnpO5I2uTtWghsC7Xv4mENcGVYbyiu9jI+DwEabIiDXiXWqfoMt
75q9fIpd19tBWjxVpNxHUHzzIU73U/4+IzDiCoZ6vr0vbynz8ka+PmT38gj/k31E
JE4qx2sVxZsnykglrnyDl8M/ATHOL7XSH4xV9HSJUw5IRUaNeZSKrhE05COniVh+
2yoN5T2dSlfLFddYey64pHNYC9x0UPvLMb8oQE9uYiRKDSiw146BePa8w+rI5cWh
EhWm47Zfbn3uZz9NqONNWMOaVN6htuvnUOvPDzaA93I7LIkq9d+JfOCBHt9fVlMx
F6SYSGHQtYJthQv1EzRDsMCCPVpLNC5Nnu9Wy7Nn3BYAZsP3AACGKSSKUeRBOs/e
ykA1yWrkHjScNpeT07sCvdhGh51813QjMJMdLoew0oaKlSqZGPOmGe0c+akMWaZA
/k1seN58X5+27QLIZoN51z2324T5JPEF+9RZOW0Ym6XSD7t4lmrI6Pg5ASTHQcbq
YToRNxG7aUsGrHuOuAKMChISScirV8+Xjg1SzqgFZC+Vseh68P4iM10TYS227MN4
DWVUE8ON6K5Uy3GRIynj//riRxaIm6F4y4ZLXJQrRbvdfmuHygHKKw6MKM5pL8ge
qesoPqKavhO7nMiBL8+RBUql7c2jt7fIE9Ow57UgiL+JoNBkveZIIOBLVK92EKp3
tQAkvsyk7jkXwqltJCPiAj6aelMq/1gGYpw2fC4IGDp4eFc8s/FKrLb/cITEZGmB
7NaZGnLN9L3Uddfot0uu9qalvBYyh0lcnhpNbqbTMfEms/6Ck7wGTiNwpZO2t62B
y/TcX2+ncdnWZFlWKOsMOgh4pq50tPa2rjBASDKlTib7l6k0X62Rpa4Vk2mREcmo
9fNcL+Pqy8R5440NfqLDqruej9SRoyScMCqAFE5f8wxnIMo4gedNBMuVpjRAqv+2
cZSmI8ZwEjkaSno+4iIg+8M+izJtkq3uucy8ZAN8pzhb0k6tYe5v/0Cdmac9E24N
AkyRgSw52qxW4SjQ9G5uKthsQRpLyy6BVqifjyrKsAszbMUyzd+BAC8PpY8wI7Rs
P3UctKL6LpAhubCXGAuRSIc3CVQIYPkcdf1iQKsXhuHxXL9IgRsdJ+cZcE4KHcGo
4z4sjKYuNofguYmopRAyycZiabcLDNeT4Ttsg4jr+gGrA2gneeRzJvI7IkJw5+bL
2HFSty+fs1xPnOzRbRnH6/FrSk/+VyT1b1hZLijn5JAvrNzhP9ZKYVf2ruVSzW1d
auGotJvpFmgtX+SSHdpsfAJkUaoDg45BNszRbPGd7J3NpG6czjJSJxl6vUhZNc2o
ASleQnZjGF1BTVNS0h3aJjZPzLbCmWZLjHVKK+Vza7tawPi2M5+vOgupurF2TNGH
CyjrWBRtrSwfVAzJA5N0twBLpGKJS/t33ixr8zKeY0pSuELBr4+SXj1IYa+eYcC6
y7t73e48BsqFjzSDXOfv6pQyHryyt/sSAxQ0x8V3Nt7g/2rdmlFkNpx+0ylI3lMw
Cgt3U/INtSTGkdrny5sz0P5zhs7QZKaNaJ6mUYTuMLeJKVMLjs4MJel+5xjW5WCR
U3jWUO8xZLMb+0Jr0vILkTU3QTcTKkYwSEuwsmS/DKh2LfPLDsTZxu9d2HB9Hk/N
0/09uB+C1QDkwfP62BjdHQE0b2HYXOV3AJkWa0Lb7xETHfvD/0y1nvPiWysFeGby
FWotL5ZglUgSj3LC1ZCh83hnpy9xrPdz8EJL+mvSLzmPw/eZEzfrD91AAON79lIQ
OmEeo1oJqv7AbyiQwftP+KgErZG6Xb+W+NmTlopmhW5P2ZDYNuPRV7Lp/+f6E6PL
Pc1Lq3a1D1ipA1j80tPRkKDGnBKJE8MYbXTpZesBSbptrD+6yJEyadcF/vNYCaYM
QNhD9sDPRbsmu4Fq+2ldTDWu0wFAECEwFBik+E3Mbn7huyo48mu9Z5AimXpTpTdO
mC+zOaf0Pr4zNJYPYCx25PCuMjBXuBOzHcN16iOUyGMCv679paL6CixsyokG0rTu
08DGPy9tTxIM1ZqGk1zj0xqqMYoPHDhuwJc66jK6fe21dnTaghCy9S8bcntZaJri
er4cinxUEqYvwhhe0qn9POmnfol3ALsxtnQl8YUODgmJ/V8u+6QLSMYbDZps91vS
plo40AjxKChqP7ocmHeSMVudkULmQfsEk90BirINo2tkvApkqfRAzAq+Il6ZoZkx
lLExa4ss4OSY60/Kw/o+lXUMAjc9guRA9ozJjPokjllRRZyvWG6dVEPDWoZBOaO0
LQVCs54DKnfTELNzD6KLj7QDBG5A5zvfvLwxlVl8llVq82DnRq+dirhtWS+XE37x
X9PGKuwZvrHvdLjjomIR4kHLQYrVUcrOEBK6nTN9IwNMkiKdElMwCtgL8VU55cPE
dUYVZOYW98lswIblqtGzMBFuftIetQWISq3TVQrIE50D9hH6hGmxypW4eqzG4cPh
iTnytjy4Kupuh9DttI7PDHcz7UCofclFeRIj3pnvxQdT1xwwjxhlt+632qLCpUKf
K6LSCShXoIoXtCasSUg2OLE7rqslfjY7Tf+Zk7dM/cvuKT3slhd3oyFm8PcXgWvQ
LVsKbblCZH/pRqj/AgMM9K6ALYnKhoml8WLdONFtO5HwM00bzqPS+CBvQ4S7Du0q
c8LuaM5z7J9/dOJOuF3EaXF55ZTGC8JWR4uYKgAEg4KtzG5CFaM2tIm0043qYmEa
mOjUg0IlH9HPJ3QKOF8bCVVFww75WsEK9f2IJQAB8DG/7QtX5dtbrbafkb3hkdJs
oFE2ZteyqvJKv/zgvUxkB9nV6sIEnbvA8bsGgBcnjY2I6a7DeTCQT9tCHVV/S2u8
86GS9sVGwaUiLYAHiEg4FdtroH/iecb/xOROlA4O6vIDP8UMluNIbAPxESgCRbNl
Mfl263mLhZ5hYVyfTiS54D3QdINqYx/khmQY7s0u2NM/JlSHMvmFfvPuuWEmWVRh
QpNU68qJzNDDIm1YpWG+bqw+ngU1+pt+HerwWFE3LS8RjLQ8y2jJJXWlb7Lccwb8
RKdbYoG86XeWYgKyMWrvyypcU/xHdiLc3w7jgUpP1EHeYTkCrn6UP/XJwMb3Ns3J
4vUNUrEa3p5EWIX9LICeOT6U2GdiVUzMkFvFHcHntDDj7QgfcWSi0lk3e7Mpr89t
g8Vkl+D+Nnv2kTSJB+NCVxIy1N1iaB89OLCLrKLtN3Zf7XlmMm2MwlPJkMWxapeS
CaqFK3sd4kzzHBxTez+65PUXR0CbNEcxPCz7k/uC6qtxW8JIZt2z1If5jyJk4dyp
EZUhKfdg1LzVOGN4XDVsdgdTqDETmG1rcEHeA+6Eid5uEcKCtie95PbyqQeAtjkn
RQu6+Vsg1pQ82RamvJYh5sBjHtYGJrHcwHJ778Xhra4w7By/61R3OZT9hxG29rP+
HACWnREEmGDMI4FQjpVAtf8BBbbecpvoX+FyxAVtDMTcjHm7tVdrdo577vlDMWTf
Y7StVAR/AjRT0PVXNrNkamOU161Ihumln6Rt0Sgk4IIBPiYkZjiann03t4yQBUQV
X4kP3bZ/BsEMSf2cK7C9wHqQBoYHo0CUMIJKvrYbe57Bj/cSLniL+AjUOZbzwrBl
Z9xWrAgNTcLCZ/OfN4WPUfbfnLkWeUjr+6EaQxifRuXGJe+8dbao5bLrMPGQsh3S
EPNESKkW3HOU52AzEUxO1CW31RIb28j8Zm2u/RXu48HQQd9QQJONFotjraeDUhGq
p3MOC/Nzg4fWsUjFMzDwv5jEomRiKroM5sMHIzXAd3+GUQifLOhoeJEEaCNDaK+e
DQVOqlSO82ZOg0BKIB/EQHJwaf7P+Mi2mqV2Rqj7+d2FDnsZj9+NCRs/Fjg4YZwi
rip79nMLnMPNxNJmH4oo23rbGC8ivbHHyq94ZwMg4ftDOBgRT5xJK/7RB+XuKvBv
D6ZLNRs+CapDAnfyWARw6kGZLWBQUXEqcg1PiDZewialNdQ6vmLo9FncDLab5P2I
/i3y/8jSIo5VpB58nBNwmxuzMdbAuPxNXfZVmtyv9w8kiHQuUxpVDpiOdj+GmD4I
PqSWjCaWcr39WdVbWhItTRvXRhRjio1yYVJw7wcRo+24Wy7gTvnBb6uq6m1CAg5Y
0VA46vbLkpXhacvl2ysS6nGfRwaTMlCPJ4WESOxIeLfocNxQwJLMQGUaX4jgo4dQ
saIGnsjf9bW1vmwmeLAPYIEhkRAXAlaCBvEOgbrqvhQRL5h3v9//Ym6u1rYP0jvN
6TIYHotisTnAswpTyNVHJSe91r1Yptm0B0bp36PFrIJwuVgiE3gCINhImiQa3qaA
MpmZW0Tj+g9Y9+wOxSC+2pDBtLQeo6YtJg1Mt+WMyOmQ6e+/euvgA2xDrofZl3ND
pwOzbdgxy0qzYVEfuBPsoSdNbNAWiAYl5Le2rROe4GoL6NY64HwfChWUONl0yYnJ
hTPcbrPao6ksd5Tu6IuMGjNuL3Jx8JcpGaxLuWjNZ/RYeHA6nkccJD5pdDZ0+erQ
3qIoMu3w73p6lZcRztmtMxC97YdhfwD9zEXUthTGXqgL+0jo0+Hq/3miMX/A6rye
oXCItoqDr08Em9xMLk7s5+I2JkeszVNt+b7ebOTWVlVo1yQBi6c73lQoG5et7Qg7
XtK/qkmzk9vyb3EDkOzNqXYOmJws0AA8XD97Y0owifL5Qmgx72+xd7bdyrLTQMf4
7Zy1+srCed1lmJgel1gnzbHVweWCfVW5O+lz9JP+aKc7F6BA6tpVNv4lvY4HInqw
skGnuwfPGdjOppRKVpAqqLDzuGdfFXTD/njV+8xtNOWTOWBkvwOdO9GxlHEp6XbA
Hu57dFRrxTcsNzY2sW6qoZBqH03wFXoRrLQDhIqu5TDrLKRZKe7/kFpNM4Iixpy6
JyHbnpQeZYnbzOyA75iIQoUJSYr+kYMRedQp2+J4/4NpW3i7/mCzYtdbXemmeaDF
62Z9kySDpl0u82MIJK0127LtDDkTSC8LDJUb21WEhbbhvlmoxi5FV9DZQaHws33p
1bzGnF+MCRRoJE59gbt+ffK1ORo5wXm8sARUI3sS2RmEjuIUnna68cWCSqxl3ZeV
ywdjatoOB48blQyHpBLdM3yU39XbQ4juNxnGZMVwdj2O4vTf3SUVDkETUetfOQ9Z
sRMfILQGp2hkpdIsSU0pLZZPWjmb+PfZe+kRfdjGbiYACvN/j/aSEbI5ERXrKeW5
qlYmgXttfQB1yH1DHupXNOhPH7K/3ORMeoWv+/M4ZIAO8QlYmijz6DI5PoHgtQCW
d6RwyZfM79eD+q+KwAZ2MtxK/12mOFx456Dg0ix2II9DZLxj23ierdBzimk3dgD3
AT4N67qtetSkN08xygDtGsW6PZDnOx9OvbWTAqZk3ZODDmlB6ZSkUJxh9mIGjGdr
If92mZMQxxzgitH0Y+Xqr6HeisySlKYSuL0Ju/AFRYz+GRyir91rDLG7AWwhbRi9
TsCQ8DpEPN0yZrxA2jSFEEpvFkEf7dyINabxRWL3470l5xW9woHsGxtHWd9S8ZUS
qVKy84mM3Tb8zZ/DEvTO5S1xEGPz/SeuvUlQww4xOWzf2wJO795wWKU5WSCm8fK6
/3XeeawlZgCadRC5PFljvpUjjjaus5ZoDDUsGuRSZWDL+y5sWQc1z0sP3cDtgZwe
K4iOmOEfqhasQzJDp6mkAea5UZ/f3b18xJc4KUAMIGu30Aj4b+5p0ASgtzos+gPF
rv6QOIdZs2VO9tngfZrG6PrXsICOKXfM+VBfA7scX2AxeiY+BADvXZQuZLp9XBo8
eR5ASXUL/u+NgnQb4JFeuVQxq56VbRJFduihyRIOFtY4mnkN+XZg6BjAP6k00YhO
onTueNclGV3iQxem6gboZg/BPOn6U/PQKI11plSrADXuAHB6qt8fbu1QWzEQRB5I
9UxmHKsjbC9/TJ+BRKAGf4TwnEktUAyLu2jV67udDKfCgYeB3w9y9QLCGMD5gFvU
k7jpp/J9Lizp+JkVIwtP1ngABu3TSc9dGLRykmeGNVC3gYUqaByqHKeyYojt7UIq
V4MoVCRbgIdBMAa9qdPQnlgtXzo1lpx7YdrjY4/5M3z/CcsQUE7Ac4jrkPQ17j5T
vOJ8T8uKxCNUmJXGKPb+R8ivu4H+ifplK3ISkP+9iaPG5qvaqy59wh8Ottxskyk2
sx8/H8Eh19pwcAGZtJIz4hzohGvJieAeXd8GkHtGxyiPVRPndTiLNO9ArqkO0uRr
WxGaIYAH7I8oo+rVrUtiv/xJwtbd11jjJfGlgn93MRSmvLmmm52n04vrH6X3Fwih
YsZSaUMXGVADrqqJL1b0b7rHJw3ZYZjk0MHnodLNVti/jIaTcEcD1Q+zrNjl/Yx0
UIPvwTYkm6MeE/sLvMchkuUIDT+ldGpmsZCrAykXFON/k+p6mAOEsBoPAo2RbUzZ
MKqvUXwF81ccv28eker96CCcNi1HaLM4fOhLLM/649CeQpgRNKyPNScv9Vtxe8aC
BQSacKD2lKz/Ff9uH5e2q3kQQov9RfrxtqMua6/dXXgJO8JzP5QRYX2BVJX4029n
V875BIdx3w0AgT/UFisDDYMdZIWANx4bbJrPld7UljyQO9dIVI9FvRyGWe2D/5n3
9ccPyGaEGMuwILLRfw699eTIQOgDwf6MMcj2DCAPaVfSImr3aY0vj3u1rQ3pHfcd
AwWh2Ql1TO1yANInElgwJ7CrhyeNuE8Qb7Fx+VS9FiPJkZ/AVP3aaAg4PwD+m1zh
3BJRCoDtMG1fc0UkF6myNghbt7sc0EY/ncJnD981rMLv1KEnLhy9Xxl6Ec9YeOij
SglG2mFfTfCoA2G/dhMuqiXExFbMD0rPHcKyygV9rTUul0dkmG+mpexpGAtEFlbN
x4dijdXrXApU8HLGcXGcpSNgxrXC7TFqfhg/1/iLTo/QULS5SWjn2CTmXjDVTV1V
IC7U+lmslckBUxIgioRGpLI6NrO1NOeFEpoU3r6/t0jNO1WSmMb7QQdiEWwZ6hC2
cTjp3ZuaaiEdorrwJug9rR/bLQY2WdX36bS0SPVEDSeXCxFbJa9MtMDQcgStVq72
MS7Q267n+j0cpjJLz3Y69cpBaERv5FgrTSycIbX6S22ixTYzQwA88/VeqW9NTx3A
KZUgviGF29uYyFa+m9muunzLKmWWrq8H4g38QwmpeOwgJO+9FZ8jBCDZvgB18+Ct
PXRuqtumtnVkMEmk1UWytlB2YNyNFliyJPi1cSU+zGCbTCRCij7p5wUPd5eaXOhU
71ZwQX5g17PGOmfJSpDs/qCFSFtevCt5Xp3hZaFEJ8HzLaV39bBhfg4+QfgBou5U
LkJj8ZcwAdHJHr/5kgUVsMDKB6sQQnerGEKu+L7QU1RgQyWolgo/duwuGxcngvof
v61/H8eSK7sxnbHepy7Sz/vKxX6DaufH7CzvM20I7plGNVdnP+wr9Z9qx3mIvWe2
eOvKrWz1Map9qlLQQ29yGjF3t1GdjbbnShZDHn5k/ofp+KNRQO4TGK0NTr6yC1gO
AAiRopoSNQGH4MfIU6+xKyFIPa0f1yPdIjnwlx99mN1lVDBbIO24qw0Pn5xKe3v7
/jRzMwar+P00f23Fnj7raK4Ywp5V2c62rUg4QtUSPy+wX4UvRnJwZ3Suez2uAy1i
Z0HuieQ9TNaw7HqMqrxwFWjgBuzrxXa+WXTlzA4MVfXQfn7xvhe2IJzEkmlY9z7u
2Kfos9+8+FXHWKFAfOYotnHiKZBT5/s3BVOlcT+sR/HFaKZMg3FimBoqzlRiVNba
nQUW2WosFLOnvR7NXCJ3eZCXdZ5Uk+1U74lSxHSTHiOaXTchmPQm/4sNZ8A3LFDc
yFfcgSvVskyl6ae0O8W4FDMw3bUojaUscMddbAkZR+WYslM+RWdEhAU5VAg+3/Qv
aJ8KCNEO/OlyZjw87w9sOSbcsW3RANp4LwxTiHt5EP/W6LpS6BK4Dkm2HLmW8qUC
clYZMTXE5INqFEzaJ5xKw/ebsRYtpsOVNVia+IVW5UZQbKqyfYnoTJ/dDT9Jcgon
dUscPD9HZol/8mIYUDNwMVhzAJuhSp8nTwbZc7KlRQ8ndx2oxQmimbSTsx+R7tty
s3QVJVQqwjUZt3HQR8mHPlRIdXf8X+ijOcaAKNwmZDUes4ufMX14fP+ue97b8Ppw
yRs/Pq2mMZ13cQKp50cPZSwWwfs45PetnRzJL8btNQ7m1+1i71CkeirH1MotJy+F
Ep5ZXXIq3Fg4adXktkxw8YfC9KjFMkmblR8sEnmUN++CaTuU/CkJ+a0iLrQD7BYF
Ki6F2Qrw/5d42g7ouXB68ZWU/7FmqU8s+i05g+ZLxYJuZ8KiO705eJs6pozWehqD
J3ymnEykgAqdQjW+Sh2pEIGk3t0jEC/9EjhsfwWntT6FvSUzVQe7Gcr8OlnSjFbA
oaY/9e/nYFJPOWJrC0fQJqX56Sv4qOTgngeT0JNxbMfNKL4oxv9vcIrS48va5z0M
A5f7FkAdmzxqXpu2Hm+uIjfdATuDcQ4HnEwMDoE6DM+uf+T5gQt6Zd2xIsgwd60v
vaMEv1ZyZnow3OLEV5wTdLMlG5m5fBIoWPdb05yDEFF3G5yvTjBaCXtnhdc2ye8p
CduEaeSoahPsvXmojD55KLp1Xk7I/tFlPmNdm//pyyMBmJ7pWEEpmiRJ5gEvj+Jy
SHK/jOrlUNFXameZwrKZkNzo6ayJCShQBVXDDxInDnD+u5/0z7r7SWB4y1Py+0S5
zt7cmOVyE88hiSMuRvlR7EGu03fZ4NuxMvXNt4u+xfXHlxXxdD4UOqOCrq/TpNip
kEk1I5USqeOMnZJeK6y3JSfoLxHHWkjfN45W/YLOnYZq95cEEm3ofovCdEJy2Mv5
Dxa6x8Ctj9PMamVg6wDvqZU+niFjViaf/GsUPLTipLoR7eErutOex7AWgczGLh7N
t/gt9pquhx/I/4EXlsL1zUWVi5Q0Im4zNQmhCQ1HxbY5tJZtmeV8lrqxj2bh5ZTL
FaOrYJkgsrQSR5kVG+cALOHSPEnQ0dd2jCib0gZ/eB+O7ykP094v/YzKDRu/Jttt
q6RQXUMG+tYUyv9noxD/g5XRbHZa1z0S9Y261DrcsqtvAzB6yYOidATzItPbm96p
VOsHZl8OmZvxQYbXZTeOhaXx8VXNpscYzYWOq9MmqJKus9DAIRpj5+hymtjsjnmZ
oDHE1CoLuKATo/lZCT3/UKROYq1hDhoXDWC8cA134MXJFq3unTWygb0q95M2s2AA
FWIUJWY4VJMqI6sDtuXrW6MynGQKDtn+8HK3uP5vBkZHMpL8vECazcoFSTb3IX+C
oQuSXnEzi9XpRi6q9Z4f/AucSknE+ge+o2+aSEctpQ+RQrv41hxV0fiuS5VohdHH
7Ahftj9Hc0JlGXaUhmYyeVGs2kvo5OwYUTshx3Hn+tRJsDzRfboo+yGQn8WCaL5W
zu6DDm6pHKQF1TdfBppmx6HfPFMFG4nbLfpkZQ1XGNM48KEaKhUZdPNm4NZEgG8Z
tZIcx9VvkU9D9HK1JD0yJafXfqAL7zXN3riCntx2NMp+XSa4ZQRX7obSYApBuBDz
h/3Xib7mqkwaRP9mstkb9iF/Pcgx35SH6fYc5hUa1wC7LXsD9sHOQBKmF5SZyts3
UkovL3oloaOsqDZcYkD3z5uf1ccp8W4RPVnBZZ8an9tc3btexm95z7N+xZxqztdU
UoOsOj+m7brui2LEqWhSWwoPk/UnwnwxZWwJ+EGc0sqVCEZFHW1CnTGNM7b3yH+J
qVS/tyib4ZvkZo9xDrvVg4mMzEdanKJrBFY5GeDQ3sGVDu3OEcY5Ji1pokqH0UmT
H/1EwKeaM3xW8BCYgFGlTF8gyPfuCexrsCRvJcFtTX8+D540JIKNHuQ9tOarBU7K
visILo0LDE04+OataOBqRJLbik3NmZ/71qKtBgZcJn36czkmOaxQ5R/HFKK3yNUs
rKaekAqASO4yfq9PWK08up0EAsc8qF1tySrJlcdlWT2eyiXncOF1/zwKYPvJSaHs
LhwRtmu/g//HL032609R4ZNUY9K64ObM1/sTnwVDJvgjBFomXrC9wbnKZJD0XoXA
ihdgrg2J2UhycFdP+bG71/3ayUrECAQoYo/p/4f/qdo9rwueSqfC5AKvWT2MfJjt
Gxi+ZiuexlaDwMFN6bia5dolhSHSh9wc25Gy6+EJVp+gNtTQXsx2f//LmSF24XeE
tJ5D+3hFpJZtipebJvCzbC54smcZNybL2PLIsFLSf75aXxYxynY5n3c+oeUQqVEK
NNTQIzwd1sLQHW0cUUpqWkT9vRp1WdVrroEpSdMW7mQzpkE34teafNt1XuvmWctu
vDaxSQIRJECg3AeWB8I/ADi7zcpMQZ94YnfUDXyi2gZ85dNx4TYQMHmoQQ0WiJuW
Hhn2ub4ytxOBVUQG25qT5jv4bMx6hQPrLnueX8rsvYrL0qAWwzxxGarA/ZkiIW1m
i/9bLUqU2y+qmJZ6FHvVDBmBvk7URRuxz3JRCtwPHf0NJF/bxbY6xJR1uOI1xBh6
EBe+Bndvms3hlrjjCfzYkWlsQnLIisEi5Sz8TmqcQous5P6kpX0HtZyrRY+NsEzI
1pcfLK1J4Zrl/NIC2W0u/XORUQalBBQ5Um3TxAaNBYecmGgre43sCOVVkLgnMZ6h
0xELqsP/hNdflfqldqZo57QCtSISrWbh5OfxZnMCTGB4rRGAd6R331AYF56LiNAd
AGf7BqVQWThf03FjgWZXAnT2QK+wbVOMu4Z8B+QqC6YfcOkp+fU2fLP33pgUuXTs
sKZrGVPbo6mTBqxYTS5i1C9JMqYxLS1TrEuX8+QK0q9kSZLBeM0WYk0z0foiRMiL
qypdPVygTqp0Aq7gAHomkzFse4FUecwc37+VJAOFWtRa6A10MSahw7JBVrQ6HVh4
BrB83GkO5DtzzBQ5j3NNOYJBt4TaRP4jUjIr9AWL01M4AsAqO4UHo9dm1V3/QHaP
59RCBR1hzNbkBjTU+9IU3QlfjI+zy7tRTAn5u/Ptfkq5RTtXVcmaYxu5Lq7NZr4r
vctd+2X4CmAxt8marQ+Hr348SkbpTvLRZnmAz/QVegeRvnUPXgnmSmgqH4ZgDwSw
p9S+J7WYF95a2Zk9dW3RXxEEq7wwVyDFtetde5Swfw/eETDYCqzOTLejehApudrI
CNRTSV3z+1cFOWVuKDAph2oqVDBRHKvRFpfgtmGj06hMSfKSDCSaKzKt4ms1H6kp
l45CFJ4IBkfj+d94K74BWrf7GheYkapp0wDknfHmcZw/aBL4jGj+njjPGGLj7tAL
gmj5msi4Qet8k40m36akfll5S4NxW8xe30YsIbaOjd72yGnJDRmF3SXl7r5Dw6qW
bscemgbrnkuCcZP3BGXBVESxg9cgZiISCLSuRPhwXaMS5sXimPcFvedsj1FTIhAU
rA3Yaj5gyu6Wy0rZ8Gdh1cf8UwOCtyAzctnrbftXIK3qY/098ykaOya5IOReHAHU
KGZCP6mtviFbYcq9fXWOfXmOYOaS3IKRlb3fWVqFhbxRHx9mHuAiw2P+JouUv9D1
h8tgj7K3JflAPYUlAGRMDHtKIe0mk8hVimh9FRZquUOgS+0lmFP3RYccrOdrGWtL
ojP9z4RKzbGCytTSvenPzvOO8d9nL4yVFaePozo4oWgw03HTRcBtrgmX14feFPnp
xzHBy3EEQlmU7qYltv8fkMpR+GxN0CxaOQjFrHJy5XdCfIelUcr4pNqbIAjhVtbb
Xud4FB94ATOwkhok6GhjKkCawsIv8QMKsVxxWwC1c/6jThp6Xe4vAEpjGjKY3Nse
FwKmtaM31gs4Syfdr8NsVs7vQcLZ8aeybYfRQ7CQHkf0eo5Uz4OAu+qdkiAUVN1o
DocY+i6PJXAO9yL2c43MXhdnA5cQkpqzc+vWcZ5Vi5sj+gDlOhY0DMCqtgrtZYtB
nEuLVwwsF8kuGg4r3YR6P6l42FFArMK38WSad7p44Y93gyDnvAed/Cwn551Yhmma
SeYxKmb8zS9aeyDgCx4TD3SmUhzf7BLo9Ji2Tyx2MXIEans7bjM6tlTxdFppHkha
ygJ1guiHmoo0LhT2OF7B800Q4rFFIAwBKSzU79Gd+9Wp/C2kMM/X5RrdYkFY5KI+
UJBLQw5LzU3H3H32K7LvIfZhpWgWT4ITri06PML8ZPkU1JoAeShCV3KIS1F2vgMM
jWyGSfljLu+bWFWtB375P2LL7AwXC2IrW2IQmXKV6Nu9RhJgMCqCrN8LEbia3bt2
ttqAfI99938lw4v6Qa87vUPznKTpE+gzBh+7ROjcZYglGl3jSb46/zYYnvhIVnK5
cXBo1hJ9naenQn/8ej7oZLmsNBf2Hwp6/dOkTmj9EuXs/4Mb8GEOV/swjHSAV6r6
WAHMKg/12nyIITt1yZ3BH0NWI98xnIcdUyPLm3UYY4005Za+m/6Oj7lvMPBsYeo7
uo1iIFh0Q3/gI+vlHoQrvqEQ78xFmJC4S9IoPBAFndnDwyL0/9kUFxG/XbcY/QGd
MPVMqbzpUWrXsI6hZJkBVX8ystwEqfghQeRHJLu7VpDIcJMb47xM+Btu+d53+Rg9
h2lH/XLtbX1Jw5AKtdlpa0/qA1oyEXNf4Y5w+ZsAOOqoYsBxgEPkXHI4G50WCjOP
QWYEZubhlCRFFLuDBnKwzoAyq/cy+WSeYqjb8+til91bgAmgTFoDtI0QTrWwg1pF
ScVdn+XHN5AFz5WxfMTL8AeWJb/V0paX0sX5TLhJ+8RaCXa68dOEja34zNaLifMS
t+ubfBuvEoDT9YgzJ9DiVATefh/FJiAIIeUx+mRrDGkCJ77ZBJcjGqqueoVYlIQB
UHOQfB9sxZGamMuzYFbzjVzzzIXHucFXHiB35W2ILLc1o/e5TLGmYC17L+DniOQ5
vZrWfdsrHgIkgCdfMIqYor7YwvkdGOzRu1MUP/NFOel+uysJBQp05ppoVHLt5nJj
8jCchss/agPHoMaY4ot37FCg1w0BxVcHmtuVNFaNQfYYr+Zt0Y8oKl4qapq0KVPt
d867DBKFtc5ovSjfno1RudlTR1tYKBDfy1Jsy4lCv7pBJnGlIqKCmxqozVPacWCs
oy2/J4bEKbzEZVPoMMvsszdB0mXNDPc+e1/swGqPBeXnmRCGhFnz1ZolHaXSzdON
YwnfYrx4eZhyS0P3IxeHhaAwtCoSzWAJWJ6oA1kK10wtb38m1s8coRIA4eBRvdrx
nhONMPy9sRqPhWckHetTZNESeIDRFvrA2lQgpAFgS4K9Trb5W5VJI0JmnEE0zy4/
3tCiSCNnHefqEQ0BQnGHM97kizOdIrL476Z0RyvuylhgN9bWc8kV33Pbh6ytuRNq
+88qs3FgKI2vNcb9ZWLV9ZsRZSxTdfm7Ux/Yfs3acANcbBc+WXziwJhC1JlmDbJ9
q1b4X50Ovk64m1uH4BepCQ9tNc8G53QnGzf6714lzVwDsopOd+EBBXsUDhrleVCy
H+Gkjl45ZMDmP/qVDIKH73KHfwSfpDO+NURuqx+6gMbpcPSD53XIe2ks6xgOGJBr
V/eU1WmBqgMXO4jtQtU9IX5gryjgtDKRV7EnLyhUduG+Uk1B9x60RDMwlSox6OoX
+oMhJYyjn4yQRxz04tEdP7By+YR4tSmDAbGI56d3PSzHlPgBSkT0RRewwVbZkpuG
syJ3Ea8r5x56MnmdCf+fhRjC5tiLwJTbVdqRCU+leijjXA+vwp7n1iPn9fy1NQGy
KzeimWm4BF0QEv0dBdr+xOIgffYCFKO1GLB9rWTakD8+nHYpFj0KVcskknm9GHMN
LZyt0LFWnOJmRRixaD0+6OnCyqVOdFW8zKoz1KBEX0SxkPTAIsze6FUFbjGdqiYE
sDuN22D+oUOV6rVbsXuZv4Skklr6kuA1q0SHhxbmz0xW6+1ybfs97mqPU7RgPho3
ZB8ntA3aJrJq41rBdVRfHw/2t6Fh42L2JpnPRAIeMwHQmNTWfc5Ju43+oRTkYrvF
c0NzasVTtojj1CJKc6sMHABenz1OFouXiyg6FRDyX978i+VFZahhUg3nmE/tCnVR
dNoCmy5FjLeVeEPX3ZLLYOte+i+c7ghThP/egJ1Wi751u/nII5xNaULaZnrZoCGX
QRhABwrkFfM2h/ITMto6frGlgitY1W28/AA8/IOg5hFW2N68uyfOzPyRl3NeVSGQ
Rvbm2CJl87yZ4sQehWD2DbnjRan3P84TwZZHqyq1+D3a9HSFaUL9jNuGAPBWBumM
ZwTm8ghNCuoHiEnGcRxqwdJ4zrJnH956oMYQB8DZbZMg3H0P4OU/7hXTERmD5vHG
LjG2sFoHuQ77SEakTW3JYV3PNV66GCrQEazmmFnU72ghBCDg60oq4QR8gbQkMKQY
Sj6NoJYg880IqXHCvCk65qfxnpNVgVx0xYhDspCdBLoO+s4SH+3Hu8UAgMtVMrKx
k07Rzx99YKTORPi0Dg0e7CvRKj9mYObFV4jIe7WbLxt7BBSbOBnDpS9iBPa10BkN
ZcBKNtbwElTrwObAtH/ePs3UbdMqm7UhUsm/XbCib2voleRkMrJF+NRP6Yg8hyb6
ka4v2ubFWPu1j/noJjGl08KZt6EBQab27oNudEzcI1ayNVcohwTZvycKpmcnG82p
dNlDVi9iBGebvUuBaL/X/ODKCMm25yPT7LgZLgzLu/gLTWsWuVxeMhNcIPs7xN5g
dGVXjQfbtv8P1VakvyGvjlhS4rwJSDxwbm+P11zm6s2kgIpZ3X45Ti/5dg7l+/qP
1OGcR04PRS6q36GnL/1R9ptOvxWdOusrHiBe1aXpIItnhYBMdEa/kHF6Fux/Iwuk
mOGChWJRX8Sf5ao+aHmamAn0epwpjmiX4apvsVTMdgEqnqi85OgA3djNQtsJqOej
gOq5VVsNjrVQihoTzbe2N+B6JVil3Gknxj7Yv9dMnOIX29d8G6bOI6Rv1qXcbnMU
nCCjqvMhok2r2p5SmEM3j+2jNmaDl0OW3z5lpqAL6ImNRkiKTK7ugrBaHqx7IrdM
MCCgwXe4hWnxcvg5TvS2+LDJNYoiJ/W6y0WmvjTGr+RMukvyrcLPd0sssZYoHHcM
5M2yQjkVVxcMIHFFi1gOFC7Pdv8CVobvcr8wEA/xqpakZt4PZ9+cN62WIUlijRzB
mGrJ51DHyNz48EGU5KUpX/z3Dh3NHLdB2fG+gjWhADTRi3Lv5mdtptk+GdkDMXL7
7sHEFzPn4m4U8oPgCVN7KxrzuOeNqXAagJAvD/neoeCwjs5jwHos+bzFMNJ/2fgx
AAtEkYpv7ZL98DNKXxSTwGCzkDSXlOyfDCEtonrwa7fMtEK00ORb82dPh29p2g8m
WeADpIIsmPrIHLzPzttAXDjODee5qiP4TIxnADIDNuJuOSD3twFn1eBRRQRlQY6O
fuxAq3cpY/sFBDdfi4BHgZNyxOyC8XAGKvC3O1VBm+XTUH6XqiR264OHoR6F7GJR
0lbvsCXXEjRbLdmps+yJjF9dHVFfCy0n023BhRpl1lulGP0lxJdrssYbKGZD46y/
r6F2S5G9qZnWFMJbtNeGLT4RZj8Adibyjc45oCuRsAocxt84jSS0EQz7fC3rIXAm
rmJkNZK2Z9CWMAjjWbfMfyeW00CTxwAqq0G3zrGKar+qoFJKFqTG5dco/LP39dx0
5ta/l7Wd6Lh9qd9umWX4EgQla52DysMCJcv9kRdODtndcicbCwxVCCZ90mdsF2LG
m2tq/Cb9IreCxKNXh45Te4SV4gXUmwIG0uEtdw3ge5HhLY1g2sEbROLaiiO/MAp0
jgcA1TAsmpO5/1IM21ijEee1zPmh+n4xqs8MDcD97r5u12lLKPzYLuzUMY3ZFuWI
B/y/QnO4hOkssks0jFc1dXnYUkKFUIIHWgQwowbSGZISZvbgXxN7ou4iW0egj3LG
hvKeKn/Ft4pIZMBj/2kBYHlBCJUpAWF4iQedFNKyM45ulmtVBJtp+C8ceOKOGi1z
uCqR4iKdZjRwwSKcgBs/30ZTz+cpYIVNCgGFFqzYcTAYQX+MzXZoLRnBBq9LGLb/
UXWfnIgr50SQM0cION3KYk56SZLd+N9+JxIFGkqMCcdLNoV7gbhAz8mQOmqqLJdV
vEQenmqTgl5czhehYCZdSuJkK8ZAPvYYXz8OPsNSFq03aojqLMENA8tC0HjtR6xu
8sX89PHZtb7jCiv4xr1jDH0ykWW6PpTW3RWS+LnBS/1svBTP8xKKD23tydoIHJMO
Eo6IRu5CbcH3KecxA/WarrN1CzP1iBiBfkQX9ETpI24tClji2ho0H69Fivnpn8/C
zL2dhFG1JM1ZMzV26TQ/bp+rOap4F+zGmL4RXyY/660Tk5veLp0/IWLA1ZWLNAUd
MvEC2psKoXkF//Lt67v5jRCzE8sl4xlh25HG6Y0CO7W6x5ljHUtdU20itsUKfISF
Ht7bkVtUgE4hjiZJ1ukz23QCBsK7BBa92dMW4G2vkVmQk8+EkO8vdjbQ8CYTRAg0
SXlR60biLv8Rsn3c7Zg+4dFhwc3pax6qLp88jg+WxqphHiHauBOAv1uOR9Rq1exA
ZBCeU3yaNWfUcw7+Q/kCgHVkLS6c2tAp328ZWFhpXxRcaheRAt9WuGt8BhM2ay+c
xnGSXmhPczgxWloe+6coa+EzJg1ruQoZsFZZpVhINxN7qyFA6VeSwzutZKkJFe1m
RRhSKK381tjjKwKEFzbK89ma4hTEuqKfiuBtFVveQnH3UP2SZHEI7Wulj2EZCmPZ
5Oc8Yk0nSGpy1BDjaas6xN0eB/V1XnXCPRqdPhwEJOM9K8ROjGTynDHQzAjNYz7S
kJIQ4fzDl6oQpMa4IRNkA1hrUcMXG379cB1QB6cREgbmzeYajg9/D6d4mNwTiduO
v54WlJhFxBzl4p4SlA73HgpiusZP/3nlioVaH5PjjmrB83au+1Gb49kwTd4jx/0B
eZh01cfZD7hTbzzHyPr1mjibWwSxumq+rx5muOAI0XEA/FlEKNsjvCU5LOH20gGK
yndZNdXRd9cRgyHiOSB6ylP6MLCdTHj94qVtu0/2s4QjRwgeOMRu6dW5w3rdbph3
myF7Ox+DykNQL6Bq2OXTMeBCTK6KN5LAGxJ/vL0biAjgm1uXjdZ2rbgnnW74TpbZ
Iisnu22lUodNni3o66iuUSr81HETizl3rvBStoVEeBYgVXZfw0ZD4qpu8fu3nHO6
U+5VdrxZbOjVkYn00BDEF78FMJnqhqSjBb5ZvECOaqaVIHmH1RcqIBUExF4Xcdio
EGEmCQ3K9pHYyFzRYGqGOk9Ujm2d4OdBXfmN2VT/61YSvotU5PXTTW5+bMkEDcxP
FHJdIBQGoH9e3gzqwsO6Mki5kWIdthUPRMrjdpoLFxEMn3PFwpQ0pNlXWwXvEtTU
SvHKMduOwR9wan1Zf5+6zsyTm8TMN6R6aYQ1PFMusTxXWx4uH077KiXtb4Tkr28d
UxxmqKa9gNrNGBAR3H2+Wh5DnVBvvXgWUwqJ34JnTdLjI45t4fsKjEgYs1DJEYFL
TQ1+Wz5j1ZSH1sDmnQRkMq6BGq2mWseyGDnJQUduSc2v0xUSOdkL3/ED+uP9nBzB
LHfykVPFzMN5htGTFEnWFxOQGabV5QZuAtfKEM1JV7NHC4W59t74AIt0tf2buJCI
yrNoMKxE1eMMvyB/TMDag0nsFNUMI/cXW2B7iRrfggZklt386R9JMTg/cwe79531
rz69OtHewGjWfC/rl8u7VhLPV4ysXOyly9Dfhk82h1MhHoBp2t0mF2gn6Ip7EO8V
/9q0oZzOlME+uUc8EQhQl6Ez8Un3EVdMiMeW9jokhiEFhUmFpWv5J7Tkelg6DGu+
BjY4Kkj0OcwOzIATFEiWIR7qAqkBABwY9neOX+QsshUx+ltFD3RkdlgbxIBNJ8RF
RSTYMn+SLQOv52+wqk5z5lBtBQMtOQcc58ZPgWKJA8Aof8ShQkhHGBrUON5bl/rx
WKqJv0yaTTAXeWlq/m6G0B9QfXGlQgZhe8giTK4eUWwpuwRPEmOTgHm7g8/B7pAU
EL68NYQ8QHeeD0rs+JWYhk33b7sJoNZIN92ztXMVKIdhuoE7z7fOEcMCpu2SNhF5
CRfO4aZVA0CtyqIE29WhBhcsReS6HYTCC5fjoaT7dqATVgzDiNTS/1QGhABRzKLr
Ku+HYCBH9jZRQwJU+XI2qRg0JhC3GiZBnRMDKJaeknkzKN2F5Xxd+EfH4FIN29K3
CuyTgO/S1cwbYEHb17I1ncsqj1KHNI+HjcHJWCWbfthwdGN5G8YDrF1YbKeQG4Fl
mj7pi4os489qn25OMdabPTLMTpe1g9vySPMcVuzooLvvAS3uGQaD7NaTe8sJJY1P
FIgE9a5/UOBxobpOZ1CMB1wOlRFG1UoZYZ8w/8jhyZ4wPMWpPJbsizWZe9FDcfOK
lUiJDtlvRVlvqOmam9Ijtu5XurjvKW/+TQp9rUcjQCB/MwhZcFlfUoo9KPBPBb+l
dwjbbOMIGxqKsJaQlFiur6PPbZaW6cp0yNVx07PZ/WfQ9tr6yhdtPcbMcRZPWq4D
4YvjWGCoBUJZnd1/2cmFDEP2JlN7mk6Z0YmoQP9ezlLcVSuVEZUW7aZR8FLVncvT
sc1ls4yfsam4RD7oI4VM0UAVE9rvmQcPOrFLxR9gjBbFXoKWlQ7+L1eOtAoA/W0c
dvnt0076IfyzLxlMYZH9bnD3LCtu7XPbRoiguK/fZyi65HkH3DMXiToFFCWyNH7o
8/+J93J/AtROn35YWnkLj6RogS4+5aFEN0SrKR/v6sNPGAt3NJ8vr5T3C9Qp/VzK
edJrim1QraqUH+B2FNQZrkioCrFFYG0Xei8UkuuP0N5WbGvv1uHkuIJN9VkPuuxj
6jL+wZ2zD59oqBqUpuseJsUEyKaIdRCMunAYZa2TGmISXWoNQxMGhPFFgPRqKyEZ
dgSeuBL24I5n30ANoNTZmMryHltHQkeJCSxLrLFpZglWmlexu/+WnnogDGz4uRWE
1u4QowuJeu7G0QOzxk07muCkO9FyrQIIod9ir2SQXxetRsGrtDhM6IJIP8ZDulQh
9w4wqaU6SFrB3YW5qUdmsNjGzRByUuc15jKlQ55c4Rqi48e0xemhCHKNgjl7oss+
IaUhmXNSB7QtJ2PyJ/dbgTWHR5Ed4SE89haiuxSoeEvkN0ufY8OuqPQ64Eyh5Ggn
ax8U6o6va8yZhapX4c8nNvo1ZdzrFxUgvgYDPNN0tZWhx25pn1cZkJIWH1JjZl/x
oknuJOkmeNZeHFn+vAfEWDqSfi8SgA8sVHJ2YF9bemlksYnBQZW78uJP649hgn7H
Phbs/ua2TbSp9IrnvICQPDXMdqKM1rYGQkDoUI5iGiZ72aPs8aj2qW8ymxgx2rFr
KSjlvAslndqQr87GpWaF+FzXjLfLoirFfZyT25s1D+bT5QzeqnZu8g4e6Cl+9zXH
UsiOkJpLF43cryJabB93Eq/8M8Pejc256cPVXDW5hT45PsURKq8uX+412ZHrOpKJ
z14tIO4E5ylJMOSlIr5C3+RiPBOdJg3T8NBAX3wkIj2cQ+O5fEpnJbQJL46Qqd6h
xG7o9CgmWQzfCPnhDj5ehqapc6GrEWR3WxHtsw99oRN9M/BakdeoQEj9C0qbpsKY
U42UqrPOqxGysYIG4TjoUZY4Oz3CIzl135sIIUGvXq+hEuXkmcDz7VyrAI2k29B+
0/Lr6toPQ4BphqXfaZfNJXUIAfj8v1f8JfpPTgOH9tyCD49N2+CQIqvKBTac7XBx
EQZtYxwiz2RVpvnm5YCYsJM2ZzB4sKa188OAlK1Dy8Pfyx/UjXTc4utQga6c7WY+
OZos3h/sU3IDugn9HETKZRW2HqFpjC3AXtp0dp2+iaHKHgSFLrjx0qgS2mtzkmRf
SyJVQatyoUudTY1QySSqJ8YVnsnb3qKR6Cffgm9qQ1EMCYppIz5mqLbxc0NbGGiD
Z/G5V8jUs5dnmmjKJ3aA4SSpOK+0/prXXhnLtLKJkXbeKXwKiGjRk2cQM6eMrmVn
2IqGLn2n5IpaXjTnVrGRbQ4J573OFU5uc91+eGGDw++iBhS/RtrD4wSH85ZbgaDY
HsTIkUjrPKiGPhPpFFW4m0mjIjt1n8py7ybDjigTj4c2XiIKXG2tCPR1/GbYWhM2
Q8EaO6XHDs3mXIYfynY03wVewk0o5FyWAFQ5vQ7a1nLy6BVaWC+mtNrP3+TtVpMc
a1MGOI2/bOjD7uxOFxUBUoAxs/b97+HoREuG5lMQ0+DVd71kFnVY0EAXKdkmd0NP
RvZbN/Q8k2GfGEvoL45IMpQ8nZwgpXqCZ+kbTX2WCGgzVqJwpdtz8qIyHQi5X6PW
jcg9fv/uUrLnXokQir8vvtO3nhrWYyJ+birpOIW1UtKS6B/jFqVFZMdXE5UGhOx1
pRgqSvdAweSJ/rMeQFpHdoyUxGNDxi4jpCqux73pbq5lo3Ygp2xvxfzxUmPw0J4q
VE/KGX1TGxsYBGQK3bp5JPEEcID2xM8Yv5KoTaDIHXMQB0w0JLabhccoP0Pp/1Zn
3x1nz1GL4+aRpinoP3je4r6btuUIa+hYLmcu9X4Xnn6U5NVVUnWIO8AhRzHL6a4i
TLUMkU5ivewEqczBxl4XVwoOJaIzsc6VW6wvyq8RMKDIEnQlJx++py1pkOd0B7Cm
X4TgdOQ/S/tX7YNwZ+kvqokYhTMmD+I2bg3K/fDZRoyENJeoWNq4IFa0p9P25lo1
hdMrim5ghk1fOA6ec9n1eChe9anQm3Cocby2QWc4pDnAXNZFrrvoZbh5Zz/5Uhzw
EwUTyCn76lvFB0tW8CD2wfZo5KOB/J1/vXI3v7kcEGDh9tvylxaLn8+OdnHjjKh2
saHOJX47J0S7FWaLWCloRXqds+5EGl2VdakwZ/wmtNKotnF+ePi8FsGxP+Ms0tF0
tHIrVgWi562LHH+3PtrzIq3G1fxqQUVux+hO3a2zJYOSpMIabuGnx6APasT9x4xI
wW6ga7j5nZeaGzKjpKF5z5ZmqgSYaQBRt38av1ESJ5bz4v8XG6FrmYNYjrkolym3
33/J2LOiUOCbhzv93hrlQkzT+74PGziDjNyinF2bDDZcrd2TCbD586wo76LAqzT9
Hz1nGdJAkWx9EqDgHqXtPcmR8+QvvWwqTUHr7AIuLo3bH5hpXXL/Jm/ygp5gLoN7
buaQ9Nhe9HCJ8/M0TvyRpMCzsothZD2HH+WJ43cUTmOSvp+xAMV0wG5uXtwxId5v
dWA+mwrmgOt2Jjm5L/kxC6K4vjNU+uktwh2OyJLUNZdo0CLPEn5vgqwEOmQvnTT/
a/wl+aUe47TMyZyDTQ7AA5RwZdpvbh9yDCkhaCdIKv/VXiHRUpCM15L3txqsYItj
XCvaN62TjIfnsMb77ZQ8jdLmpCPZk8cYPYgzW6dNYB0hFEc0Ihx8GW6jXcG3/2FD
tW7olB7AlPpirDc/HBZREfvCdFrXhC3A5IhPA/49YIspEqeWMM7T1jqUnfLdRc8i
n3j2uGpxgxWcoNAC7GJBGSzf7ZlTxLVGPLTXt8gSm2M16h3PzzppR3ttig1eABmv
tAJvRZD3g2utGiXTz3/hyLtmx3EGnRATgTIA/M1GWrJLgviyvWaMGROLmzveSGXn
vSBHoUmlt/kAf4ocJDq7yU3puqo9dr/ONk4X545JSc8JogQnzyNJd7jN9f3si2JR
T21QeVpDyeV/2VskitpN3bPoIcTcKBtNhax9/H8QyTGHdm+dfpcF5D4oyR+ajqto
5+Euh0XYLTz1L9kRjiYMv7eWp5T3zWDRI3gddmh5DNU6/nT/JoDbWj+3T7j70EVp
NCZ6eY1x4Bw23MmGM0Xy9ucAQrOXwtVAxDwSkLgmui1gD3AwiuNra1lCq8ukbXks
gwkEDBrktp6IFj53EPMH4lEfDL8lgub33FRS9yevghwZTNnFIKGehfIN5hhMNn6b
cuevg1ygshwLoMSWR6vONC/Gfdif3n0hzAITmmLnp0eEmNSiFMQJrxbR/m/gTK0c
+Hfm+xysh0Rg6AT4CBzwU1o181qQb6Ont7embS/SchC2nWEiq9hlb4XA5MVSiZ/q
rfAja0XoczQ2kPjnHNnbQl/pzg4ngMzpYNhwoQHSPBX/rLUxZFhL4gIQZx8TG/8G
7defagvM1Rn8dpDulf97Qbzjk/hUcwuH+FdHEVWiRR63PubOpew5LLqUwmuMFICw
x4lY0n0vGbzCuhRQaXAtGf5Ipo1L3ogiL77a+FJ2a0kwkRFlV7BWK5YY5sWWAyDs
lU0XshLeB9DV7JblW30zb24IAT4IGKZ5us2Q9iwQBstv07z17KfhaFufxL+s6G6A
ITEnatBNzbQvzyyoBVwyKz8/YR0U6g3QVeuZVeYUECl/Do3v6zbzqbrnqL+MfPnc
IEAx2sSyci8fAK3km/13RZiz9KhkLcvtbJgxpzVrA/wNstwqbPWoJHH/UeCBpnOz
m/O1y/K8GiZ4kQkdEEs29zaql/EGJ8YfHrsgyS1ft7LvJqMwHbzenwfsglU7k633
VEONHXX1e6SRf/epd36bQ1/fTVO7EOZchO4dAzzzbfr/d/GnRyP2W9Sj/HRJQv3q
TQ2ixHbPYGuxNdJVAWFuwM7Pay4yOGsSX0eJdHCL7TXXU4o/OIBu84ptH2DLnxWl
R5p+jaRnUBQwspiZV2zSNarqJBknOSElyb1TupYd3ScSaoq6rr4l7LvQPevvjAGu
VYql/Q+DxaWVWdk3Jf2AwnRXEJ0x3eVydcprJaDlqySU7yxgq0lN8vM8engpunzO
l7HIgJD5m7sJBFkxeUSF/uh3jItCW/disxCsUYGhhcKRYMfrZ9qfr5wys1rIZyQF
MXi3L+U8+XxZQaWz8F1ebK932ZOeM+Hdr7pz53Oc3jfHhqhzSY6UszOwgxFMpmAk
mD7wlJbrvqZEjSastfmJC2Byf3DCldPIEUAdU7MKm1zgFusse8l5xo//pkrP9fc4
OjU+QnexEKWtfh44jatRNtpFqxeglbWt6WqGKLaoWatxoShSRnPS5EURnA4Nu3E6
r4NSPsT1NZcVTBxCB/TbFSPTplt72pueON3K/jTa5Lc6hmNSwzJ274oTG4D8cVpz
Sp0H3fP8PcOY+5sjvJijDovdNjVapkNpq0XcdgbfCrCsBs79xzvjrAQcfFafyJAh
hLFHKuyBRUaRvTW2WxB0p2JA9aAbItWWiqdvVoaS4T+T/5GlA3LUBHZxzX8+vW3X
aFNj+4EVBIGkGhGoRdrrDfquhT/LdpkNdHaP/9zo6szbopcAf9N4ONkLAjkABPw3
HAraHIJc4duOhRAWTe3TYyjdJz+f5lwOQXxTYkmH/QY/27lH6aXc7OtN/PZHXm1s
Bo6XJ+23rgnSMO9YVIyv/VbbW3hZ0YPvNX+D040fZOlQAx4F6H5NuyoWijf+i4tU
Lq23hesyUxSsMXFCG24LnfFEhM0pmeR8aYU5LBX7Diac/8TaNYNNObsV8bEkmT6U
ynjxe+raMKlaKpUnlIcRwMa98SlEi9o9Xa1ULsOH/9cFvOfK6o6AdNKWK6FAFzeF
iz36mqpXYWi4KWtBpDGiEcADJHXKQYr1HPs9Qsw8R8QDNlMRXifO4IRME40pSgUS
TumOe5+5uBAL14s7rMPGuuxlWFnKKXGvuI1wjnfmbBHj8icGzeKe+gPmqwkzIsDB
TeNya6wH/vZcEMEbzbkabJOTzlet84R4xW05ebmJcC2Hj6XXc0xl9hFS0OEpE4N0
BQtARnPjV0XXwy/YJBNpXg18Ua3uAQwd+SYRIoSYn0nvtz3EnzrSGP+vhwv3s+bE
5ublG8JDzDt3UwD+OKDDIKSWT11AzKV9ODvflvhTkpYEpJK2xX97xEKRWqBDuTPY
mHjZXNkT84KrR9a5nXViDhHSV2QiB3Ft0LZobnsQdhG0EO7STf3zAIwlnymc3vpE
k9V9SKwzbvnL6/6NAFQBXWhLjAehRFdIoz9MEYu9HYEQaXil2grrhotj41wb/ofB
p35+n2FtH0LY/7BVUJOHFy/CsBjMZSPrO8cAe8xLo9BvrUctL02W4/NmPhAJj+iE
wy1fx8IY40n937SHQNIe/olfY1IQvkOqVc8g3D5tEmZRst2NboDrBCGDu0GLIBDr
bpQc7ImVMOOgAtpnvZZtTZlamgcpvP0WBSnjf/Y+2Uwb6pdGEDQc7kFg6VG8SbVC
fKdmMknUR5r1Fm+rjdpwpipw2dkvzOaK/j2UvX/WPRqd3sS9DD9UJVqNmG25+RqT
f8OJlQpvq2izytnHgXFy2a/b/7GyatOOcxfLZpQKfm9o283OwNbt9h40gUnUDVco
owUJDHtl7ejUrVuMj6pssltx8Re69VOyAwrAqfxOS7T66GjvftgeNRRu0b1AbWcS
Dnp9SxOYtSP3c94/tdwTIIqazHSxC2u6Cp9oIT9F9AkPkvOjZmvA+Y9lmkUlYvAa
xYOpepU5aUZJK3Db0LYmvVN03bxVvh0/CtWWxVPNbIzkJgr1BLNJGnhHs8k8pcxE
2pIZFVIRPEniIEQVy5BCzb2xMAdd78yE5DoK36a9XQfkwsHeE/2vCJcTinNW8izK
rOenuBjN3omNX6TBJw4h2kzeukxVHuWnTMiYS1OvG0IjQV0AU7+w7xX7zt5kRYs+
E0+x8lf8+C2OicTy1n7KiisFefdfGX1WDcDpE2zxhwZoAjjpX9WJoRg/fQnso3Wg
L8/y3m5ZFWt87wfKTyMePmfGnKJ704UlnxCs/rfYLU/43zN9CDfro8E2FxnvNvnC
+2Kin/lol2lkt6SNMr6yvDsQOJ6juTnYrMnhGtwwer7NqTVS0ypsJBYBZDjr1yVF
2qi2+RQ/UiJOUMaaITYy0BvZhyWKjYH0bTmLnXp1YepD7CO1zBpf+m4JFtEYERoh
OYhYkEvCHNdt16UvrOSzeEjXOM53/yUG/DWb40lc2y8xQ4i8rW/xjXcoX2u2CMOq
z9MFMFlokFRT7zNFb2iLZKF3mmK5VOu0IfwpR6H6Bv42dcvpVHgsW9ljeKaJU564
FMAKCiBB46dF16wYFjRMbH1yhaBy7A+jDMU/I8NBOkjVGLDt3Kf/lB9+0qZbXorz
YrWON+Z8mdb7pISlFuO+BiLK70WGwSIEALOLCmBfiGhNM1x+esU9lefF/2tg1q8K
CscEWDaQ9x61lQfDHP/aTTE9Pd+rBIH+3AcV+N4pqLrs1qczEcPMdBY3Hqe7kYRm
HbGEtfD5eyC1VjBuq2hWXUwDcF5HZFreZFQvFjeFYuB2kZPtLrKDI1QHSW8lzQjq
vR3Zvzd3rJY4GnUaAU4xMxIcaNcCIV7y1IhMx8V6zs1yTHEoWqCuk9Wi1bOqiR43
AXJLOdO3a+ipkTaOWTK418c4H/L5bJF5BiIgENM2M/tOMeq/SAHhq5fBQO3FkuD0
TuWwK7Ct6QGG0/Tr8OuXIddT9qm8SyCEkHjwEWj68T2UZfYg1k3jiyx1me9InycE
l/r9P12RGYAFy/j30QPo16wn54aB/r04dEDYyXpdxVufTtF231tJGjrVz1LMyrIY
xqH7duVijPSF9xD7KBeWacbrmIvmZz3RofXgtK6JsLIS40ElysfFrBDaF6AGDtBm
eWK6iajWaddouNa8tQy+uFvMewIhftq4A5IQOE+4BISYwZn4IB6kjV7VCo/GpXbW
g+fhE101zOdfT9hKZRxt2LR2FTTiM30BIGBgEvNLOSVfJnqpG/S93B1KDnmRZAhF
s1x8Iu8ydMj7ezefzcFtOGRukpixznxyknrQ/P0jJ4lmv3AAy5VphfRCK15B5hC9
NtIN6ZThiO+7ONU4/HkmjrgSET7R/VQhXM/GKZ67PF5okUHrTLQx7NQ9u0FGQtJU
9RCdQBvkrYNrT72fBRTn+pyrwF0vzKx5xP2G/bPngBwbfT8b+frhw7fCFG2O0NPZ
o5erHvwJHeqEIYkLzCK/OTEK6Iz62OZ9yTBSAgbDhaGnUHcxBAxW7KPXFSGDo0sg
iqnPJmS5GtZ/WJbtwsDcbUCe9P46i5pLfvus1macBkTjlWvKHLf3qGtwTYoxhXf8
jUj0q8EEPVnuqrrHILTHa/wD2J5bjO54eisKiJl2QnPknmVTxIXeQ4fB+H5Cflex
wlprMdYVA/dbHjz2mCXhebSqtq0rdBZ4Sm/HK7W4LFb1iaRpXmxXKJYuabmzVAp/
pgVE6dXQE9QaIM2zD+gxXqNF8gE8RDzWf8xFGh16Cskd+uJn+OT6nf10OQi8XplE
q2gURdEUq8806envc5jWIVuGTDi/rRxu7VjMgj5rVKRAIEdh71+wgSZDw6ayXyGS
3La5xkPSdpkKfAciHASUKrOs0MF4xDHonCvqnp+pOf8vOvyZeOdkOo/NQPi/W4OB
TtERn7H79JhemqoPrg0e8RJThN8TSn03NB+vg5mpz4NMFSndMWbusGIOjGRlS4LU
mE+Ur6aNaUtReBKXIYx0TItclFH4trgut6sH6FqzZaEgOnC8Nj+TCIdShIsxKICS
anP26008RZrl9oFbMRdjoK5KSWEYHT6HgdFhehv/Idh/D8ALTdTTsIelFwa3hGdM
D3f37PevMEoYlROosvx+Imbfl2ZSYqRMDx5WO8Co3xdHimTBCWOM79w4wqcrbfh4
JKksAOMUedYVSvuqOIVioHIIBJXaVHGReNxOtRIFvv6WB/xyRcZT+q/X5KbmFVjQ
tG6e45cBzVOKTW7nm1DGgaQZlHsLR0O1WNNtDuuD5xk8TYPCNQCN6ZY2XUR83oTg
2hO1YiAv2IKNdNaEXnJUASEnSUHOj6OtevFTNsKxkKOsVaAia3LlLFuOVTShOG1o
uG8T5JTJsGNcDkwMvLHmWWvE+PoN0Lo4tRIMfJdpdpbfE5hMGEAwDHis+lXONbyi
D2BzcQUY7SYK8NW3SXMrhE2A5mzpG/K1GfeCrzH2siDUgtT24JkbwFaXNB5pe2sI
wMSEBGPGUADh30MC+1UCA/WyDW6tiBOKysV9KT3irkub42WEQutYXPkJLdhe++KE
QjFbX1yRONVgD01Hc3s35wittv1kaOHbTz/5ddSNv41tfmzdyTE4afDlLWcUqPEa
OemY/OPQlB5jsKfQkOLPNzszmhTV6ybUiLQhV+IPdCvxVUMthPFruaiOBBKZ4nWp
wx2UJ+ax6s4qU0TRM0bt27bGXvqTibSnteWrXxzZReE6l3cC23PlTgX4acWT0bEU
/Hd9tfCI8L5KB8+YBYOfyS5WjYiCmzrxFdIyCVHQkij2bwwJM3AD35vUVhJodpRe
ojdskcyPOGJIyD/ceDTNg7+NY73OL0FxTAilqqcz7U0KcuIiEC0ay4B3zV0sgT2D
UauT3/BN/8GefjzS5TTpC/qZcF2RHTKtgFU93rs8LLS6XFb5YwWZFBmZimKSfKtV
uxMWxuKPV5HCDOmPf562J1RSUL8939kL3iWZVqX16TuX/vW1l22BCks2B3Ct31rm
l2xCsgzYwCp6wdU9I9mCR4Hm/Hebphqu0ywVUg6iTUgPlNvCQ8l5PnGobKJSwAM4
kJP8su5UVlwJz4iybFZq/1/lfrUAdCa+Zt6B6xYCf1pDH6hbAyI7x8S+maVhRPc6
vBHgCrxaDBov6qL5bj+3ILFEkd78P0C7rshr+hgiEDdaryjk+yDE7NVPlTtULSzc
MLWF39822/2PEJEkWHxPJyDx3laEbA10DE+uKwCS6YfWOM9HkHr4+LaICpGHQMmn
QoOOOe3+2eRi9FRalIvaFS3iQ/FP4Ez01u5TdLU9JVhbcDg1ty9xWlhdldkZTT/9
PBdLmU4l+Egmjmf9ZgD8Tq6QtA7TosVz3/RidhWlZh1/SzR5mEsM712jP1atpelE
dlahNLE9NQIas5BQYqGJxKl0WdKE+wAKWobQuuqSoudpeGIggouZ72ooz+Qsa5Iz
vIfhLb4QZmPt2pjMp9mrWS62MfszuAxZBZjlB5POE++PDAERCFj2sJRI24VF22hs
8rwXxtcbTSuVFpKt4GYbT8xZ7GSOa3euzcLq6nxzyGXdt84J6xBGrNy+Aa1pnya5
zI7i5iiYu+GywlG2TIJJ3MiXtWjVuJN+D+pN0VqRNvAnRBwlqt5yxYRW5NTbt6f6
upCzEcOoKVcTDUxLLVRVfBXN2aE2Dxj0noplkA9i7PC1T0lYF89tYDjjZkRGQ92N
7Vbw9pD2a/3hwLD+b/Wp6gCefRODB3l2KxUpYzC/XpCPFPGwAkejGWIFzjIKruOX
sCuAtxnrPzBYM/jNLUxixlHvxlNgFsuuyWOt4K8oIS8BqjagFJjaEzP2k/pMv1LP
thzm1r0ITHJUDaStDMUsqReVfOoZO/aXkjhuFL85+ku49iWpJzMxXzXopiMGevpY
lbtaynq+hZ8dR0UAzCtPvcaW39GehyFSo3n9Y+xKgeJQh8LG2aFeLLndHE59REB4
dytGS6huAKsNgpwqeUntII8l2atA6Yar134c3UNajlTh6rXfV2EffKbnLvrJILDo
hTWUXsntqPqaq9D7ehlJIX2mXbKPdAoCOi/R1peffiEqyh4W5LfVA1c2udX7RYIm
gzHWNP7iZyWqemgNgBTmLmaanlbVZONlEXQiWiu6yQbyAdbZ94o+u+KBy9NXrN+b
mQWXs9chD09dBOL6j4aSVd2j5FCtK5Pj1bTrDz8A8j0460P8O9nkTQE1HqZBZZ/X
JsS8Grk6UEjo46J5iGS81BBL4JDRETHg8alyKSBACydZV9fqOIhisJi4V+jlx7Y+
wF5Zx5Ev4aJzLTAXh3ZcJRGLq+CWSwGx8PD0eL8Q4Avd5pTBti6Oo1GNeC/7dhWJ
aSw7nqe3E+lxTBYPWWdqKlFJmz+YRAK1mIuX/i7AoHnULLFhtwfLaLjsnn7NPu5Q
b1YQR2qrTwxHshbgW124KqpQcD6YsBnODd49ycaoDdcXUHOo437qswnydFWreYd3
E299xxfb5/cxR890yZSpQLw10rqA/AxW2zpgWxjm2u6dJEchPCpvQgqw2yHDiL98
jE4imaJxJ/958/FmAQDbs8chvPqq9dLX9tEJ9BvfyP2DT1d4aeY4TYuB7FzS8bCW
srzcEXv5Z+BnUuJj3wYCsA4+GEzAzovgiwcCKcF87BYWwRkWnY4GSU1gsrJDfnAV
14Z4/U+fI9dwJEnrculrVsq/76eaWyfKesEGPg+dxp406qMu4KIz2cGC+oc0xfKx
uJQl81NhV1PtjvNOJswS+zUHKbDTL14O7H224L49m8YKGlqbbhQPEs7YD0Q4bSLf
9fJJT0KWoIEe3yL5DfgMrIs/uMB8t2FKZ9mXyIWf2IE8zFJwy+QTJq8Ll1je49pn
5y0AgZarBuLRVRICALboxIIEfFB58gKGh00w7P72byhlBPDqrELEFnE8geYsPaPA
ZHtWssiNlqc33tR3wdjdUqCcl+bwbx4xcaE/6OUKm7rJ+65bSn1+nV1TDocYxnp7
x3J/R0/GKjZvtKyTrcY1nSWydW1Jbq6QBsC76EFErALX+vM3yxzgIxtcdFnRhlP4
vslavN4Qk/mmTVvW4lDdEb1YZAclE5Jiek3HGfEslZrJohN5M/A/4prnUIAe1QsF
YOzu5dB2pw40iPj6kpP2Tii+Cci3zqWdnCKhLTFpfoyWhb35cOnOgf12qMQuJRZZ
ioAZpYcfLd0l883Z5kKKbef/aAhM1Vl2fw40jUsmMtFPukItMP5iUVPYjyUf2n/e
odcCyf8LzGRddt6085ueiq1QUA/S4GcYE6pXaEOEGo+DI2Lp5J2catBn93N1PZY7
/DZYkean7hnb8ucf/kkxOQmQJE+ZywkOXKMGcY+YDc6iN3ixH00sWTu4LxQZsBwA
cXIQBLefIA47pKlWQmxNCmhf/j/WRm4r5FIIU10IwMoaG3mn0oVF1nkTBhAfHEOW
CFzq7jW8nMF7a/i9vvHSWV3LGRvG/DdQQ32uHzU6vWyiezMY+fl+9RcorPJx4P68
j4uTWWb/z/6OBhHgD8ZbXb4qiJqF3pqmstr+6mbMazBlTQIB/cUb1b0ivo0a1nd+
dX1jz0psWJxVrPqGYPgTlgCfepWb1Kns3/KWBtTNRd5UDpTxxfnbLyB7atV+O+K0
M2NG0huPDGsWRQ2PTOPrYWx5CkBOzaqlTsYdhS3dhbW7vpb3JtlV1OcMKD9+zGp9
eOVeLtfHvjOF7wLjzhlhonSrrjNqPAKTENQF60OEqhHswws/tzAmY9Mc3F5zaf5h
BmRX0+dc24m4oKnBDlluBUPf3X3Klaqv1lJAaECxSRB+Grpi7OTMZbUo0ujp3MCa
E8FRNxa4vT6XwcQa+Htaeu5x9KYkfNmJv9u3l8zRaEY4cwz7svTT52MDo+vkM7kC
NNkBFvAGDfUJtzaV4XVqiraZPN3YHcxj2VvfGCovhww+iLlFfwMBRjAmcwVDoCTG
ifI/AzkLV8+zaTj/PzPFe60DIn6Ia0PqgBGN0vTk7P/LavO4yh2x9GlAgY7K+2cM
6knn1QnZkgqh3KAgNGKcjj9pHRw7qRzBj1hWEWuOa0J88JvyVG/X8i5USLd7x+/m
5yul9RdhxZpIa5gpiaoZrq7p8+/NDefn0xPdvF4Y4rGKoTNhiodK4N+WWFfIreUB
9s4XztebjT55NN1QLD+DkqzJb9rpUFmx/a5EfvO9AIzq2YLbt2XNS/dcxtxbjqWo
JIHX9ImA64Zk1Ib6kb8Pld+7vSSaolQlxVvFtCZzVcbiskVAz+pL2Bsog/xA65bT
YMRpdX/LzbHlmGC80xXpq06lHHfHWPE/aFWtRdUyxU/EqoKaGHDavuwnqas10atg
hKPOq7s9+jRkOqxRo4Yye5BnKNuAkEzL1/3y5jhs/VNQkECJoDMpjFFtke17jYwD
/nb25SDyml05lcskvj4fk5lnjj5+Bqkazuf5C1uXPyF62kFpyy6jd0yhhKIDqAZ1
QlYba2txmchHKyVeYUCIrRJmiKfKnufYgDc1xOIdqWzzy6m2yBCc22YQhXj0W6NM
zFCYeHsW8P3l6IiXB21i8Cpk31Vy7t3EAX0pQlQ9/zBioM9w5iQoP4c6OfDyFKQY
jAK441oCg02uEQ8cfq6citGgdMHpH0oRKjwc1/q6NeeoSiaNtKCsmnyZKo0cljvf
tCA6aYd+3Hit4Qum22Xbht1t71pE5v6zHBLyZ7VuDEOHXUj+gNsVarTn8Dj83/yG
4WzKuwajf+H+S0bDbCUvK3yW8GFLSamG6PXihf9BZUJpevIv63qVj8s1M6hWCBfi
qMLl8NrRm9IEXyQu5C1gM4CW2L/A31NyDhZHT3r8f1TD7p+nTmCccQDDZin0wLdU
9sPvizr8TuKg6m0Xu9N9UZYUle2ydd+eb/scyt7n2odcvggsd5F+R4iqmudshAnx
8le8YmOGxuuZPZh/cTK4SlcafRqX8waJOerDzbRI/vNi9dfIs0hmZZEy9Xo4sNVo
jFCIsweFHrgUr6ZCIT6cRBnt9ueVdiN6LjyGbj23Fa4GD19Df8VdRX55eJNmFU2n
huAYyjT9XFBbejx5wo4HT/uVwvDDnT7Sh+VMbxqndHul4FYxpa59ApTxHz86+4JB
emPVYWwyvAntI5dwZp8qJmVn84bOxdcK5geZRIJjGUWo8rgSTVpeJ6slOpjFoNfa
ZewJZ8aBFQqxQNf1cyD6wTdv1VWe6h5Nk06o9Ug+WCfuzTMkV3f3qUPHQraTM2zT
qBxaKL1BqIfqKfWZrnzGURGSiOej4uLmPjGn7+RTpj0RaMWyN7Ll3ypG4Rxiaf2l
DVMgEhopVLuGlYZcOBqJ2Kc2WDQH01PVnCaVAZmhyZ7ueFDowgGzcM//yITnOxeD
o9xf7xvT4DeeQAeadvnupGmSur3rfleOuozr8LJnDupIYni9gt4a1xSy1Lr8iuy8
W6l34TrcvmRCkWJ0le5qxVtLgOV/Drk5nsj8itVCaT1OlChFxUcQvbK/uT161TDz
zEeXzPp3Xw539VOvsaKjsA/q8nRohKJmQKY81ULIC6JP1O3d4DXCbsMTzoyyFdoz
tosq63hKe6lur7BxUqe+nwdpBy7mMiu/otVL5BYJ8cIApr9yobQuKAFXY+NejySm
ZOXw3Exrgpvd49OtnYZO12kBYR5TthnGCOA1++2HLv8QAHfEn8Pjhw2SPRIbpucO
ZSPD6dUjgecN7H26PZbobP5YDLewQP9wTuI+YLu68tpbEmSogEtU1UdNp+uSRhmX
HGIUmYMbqa06jq3nxe0p2LtzXKzFbQ/C+5TGXoSHtkL70nLe9wTLml1UPHsaKqLt
CvkO6fNf58hvXoxl0OU8kMeFCAks9akYDWWbFcyqwwMX+XV2mnXdBPl6/ZAlPed8
tzfyN0baRFLY4C7WyuG10YpT+Wug0ytZW6j2KkmQfx6ssbL5WiKxw89ChTo26NNK
KYTx/+wMmXPrwVU3Hvk61tjJRC72p5ObEEEeqFz2veE2Aaz3ha16oERR6XD45PhV
0NwL7Lc4b9mIQeXjZzSNqIOjBZquWZaANYPlscUpbVuGW+H0Id0FtfczKuCRlJQ5
njDZ6k4X3ggxI4A1PbIWKhNCel+0WCBqA9tmb9zw1dyADbR3RLVYAgAhBCldAeSr
wEC7+ZzYAstHLy7AnvDcwH3aU3Yphpr8DcGqfDV03MVneqn8DEnL8X93CrP0sHsl
ck9c0PZsmRkbQWljydTRXDTu473jUlnykNd922AJ9c46XAgsgk+cNepnCUe1luZl
TmhWZhUa3AwG26EbmFyt3INtjJAExP8nxC/jHBx3TsCE7fKKu4usvAGyqu+bFcIh
Ls+8sLvIgqckjw7YgUXHxpmolYfXR33Yyr09CFp1xhVpcLvPe4RviiztilWWbuzA
DP3Dw+Z3ncWvIZpsYXUuHfrRQbQq9vkbCeE+u/YMcg/Aztdo86whz3nycS9IxrEK
26VqWfCf1axARIfq1xd1fAiFGoImU+ZrAIc6NVirajBjNG3CEhDGSrfG7xVHc2+m
762Nko5d2UR9KrJaPQf50hZ8JNtDlU8ggUpYAMXbj5UhvBhYN0L47RhYAIpGmjkR
osMVP8POaM63S0xKjbAoSXc4gJhr8YjBEJjjiA6yroXc7ghsyi7p/68SgwYMto9l
f1QDLnC5pG1gfd2H1OAPO5847IeG/XzenCIR9Yjyu7j7bgTlfamaK4GUS0zbv3lt
fBttDWCgM570ISvTayiBtN9ljWjJ1yWu2G1e946J+uvOP5C3BprNijYgATiO5f7s
hvipNJnVB7aozrg+akpuWkaeSxQPG7km9qiE3E7J3PVoZxs6hmQxiLWBp62AR/aL
rpFiLMgJgFjolFfq1LU8sCfWCr43L04eCKnHqwI9Kupho/ks8bwlLwvKil79OUx9
W8TPl8w5oM+TMLWDe3dHM0RHYX3zdsls78SKOWwbGflLkSkaml7vy0gh++1IDjC8
4IB7I+D2yC1JyC21+D6swbYfqQ5YIp/C9clI+NZHQ/pn5JNk5xoloDXGX7zxDqi/
NIWs17l8sI7JsiHaPOQ6D9V7XF2Rbl36/5Mdh3v3c8WhZhHZG0YmtAWdPhhhLs+r
BOxOFFe3Uj+J/2rKB2yp4/OK+7DDX+p4dJz49UAsuRAYq4LwQJfE/rwxH16fIuqq
Hv+PthS6tBraymlmQdry0QMcMr7UIZL3cqPgr/8ufm40yK4lo4FdqTs7PWWGmoHJ
x4+o4Ey7vbZJwUk135dT0v9qzWfO9I8lpjut1dGeAfjzT6yN+yg/DGvhf/1Hg2oX
VgKEy9c2gvLKuYWZC5ZMg9Ui4NXfaA9Ed72bItAY6bRqmv7vOxT7T6scd08NXG3F
29+kadL5n9yQY+zWZZNG3i2aR3QJvd1zo+JY1bQ1JdJ69bnD+JXSEWsss05jY1yt
WgNXvtVayZkHmdrVt27QmGFmAtPUP/OHtR39NqjI1KUt860colDVoo/qKCSUB+gb
2JetVX2rAkUH/ExwpvETXvDyKq+WMPhpPSAMwoSo+sPMYxDmPV353Ims+ZXLeLf+
YfsSbxa6hjZBlJgY3iVgTbkeSO65pbe0APFPsS6eNxAEM1ym/DSk8zgHYJ8Vai9L
W2YX3G2avrEBZrwt+kbQPof/wO+dc8Bja2TIyLRZ2ei3UP1qyAZSyTupJwgwas/r
YZImrIRJNr9/n9nR4Z3VNK9iGIiMVWMfue4SI/BbpKjwEEJqb1pTY6M45kv6Cnvp
6o7OnJPvF/UzAxyBYLyLFvdK5RZLmp1xS1/HVoaO3BcbPCOiueSsUYBuM4CMEKDS
ufXXz4bMxVZDY2GOq5lsT5lBmmhkRPOByBY9cQrbwg4Q1FbSgQ//DwMepBDwS56L
xRRzU234nqUTzXxhXlc64kYJrRYLupSNcAGypvz49/DYs1duCS8wI8XNvKxYEtib
QrzhtObV4Z/TduoL95RMH1qXwzKfjXdmIVwMQgaO1aZeXR0NmyYy7NSQRWYXUDYU
fX1j/HXOnt404q5v8uiOrqE6wSnnKRsdF4CjCvuGF9LQrxyA/VEdntxkxF7gdqja
rXJ+1xM26FoM5239a9XAAztt8t8TVEpGzLLrW+cDjnpH6g3rA+r0zDP9I7cFzjYJ
m0qL9bzf/CO8G+Dum0DZcU9/oUc83syotKAbOet3TSI54UPGpargAopuKl1DBbal
8Po81wnMt2xeLdklv3wAG7XGbEut4d3ShOV3NwyLCGUuFWpekdO6LICHF3xoQfVJ
c+e6nshAIsFExMYu1znIaeCeLlwXtZsG7Br7qkLcYr5a3aMYfkyJdYfSo9G9CZlV
m3yhnUpMwB1AseU7x9OD8czP+h/lhvpHoPD/VebPFFo2k8s6nKsB7+UL73l3X4WI
GlsbNo7u3Xk9ydS6n8iS0ZRQMyQnr3wmCH5n6awHIqOri+Y4IPYW4nlk6KfOjraK
dbJk+k9rcbHVlOjObrivyb61CoQsN64EfCyApgrX0N+jPnOwsKGY6QmfRqeBgvmx
IxlxJ3R1rU4DKmLlrxwN72BhXbgvptCw/UpfVrgFdU0OD8FvQ4LXLCrKGJPb7FGr
hinlqhfrVrCL8BEa9RDPobrB4ISZqfob8YQYrhFSvyWDXAPWulFK8FxGkCMPukKk
o3wcphcgDH72o+G4S6JoFRnxEPx/aMiOQORTk/Nc3pNhNxOGqp70ZE350GZQa+AO
uoeQ7Exwh41PML3EvVJ08vetnLDCi/OTPhR6nj+CFvLXGhxlwcuTSCD8ezA/kmB9
J/pe8RTl2hLCnqMAQ0Rj+jx9lE9YQMZTKj2ko0/dWE61BRPP4iX7/r2aMMG4XFEE
Gr+JLukiefR3A8mzOiDu0/tX07LxQsbNQ92c7onkhirEVDJbRgHfTlaO/TJHpIdP
XCzCrAr29ukiu6BySisjsZ2rNPj3NH2ab/sw/5/YWkWh+muUJ6l1yw/Ans9ZnM43
/yBRFYKMtmobBI4IrhJORHwNeV/NQp6+qaIRgRfVSWCQhsjmCb36OOno11VqD+48
ud+8u8CLZAOeWLsxtAFHhu2q0czCiLHk8FsdPWuhH9ncRZ/Xy1blcG5tI/mRBCUI
sK4OU/xfkCL5+mnRU7CzbcJrsG8/95uzt6E8FDwSuWcgFuZnEjkOew55hhVKyuCK
sZQj6OPOpNiivhhLRVwNa15bV7YVdmdLab1r4LMF+YqBd48c1M//LA4uOa+tKsVt
g5Dopw+yYM83mxKal1R/o3KMFXCgdWZ+Yydgwlb2MdIeCSR7u3b+69NWFbbos+Vy
9mMLIhNP766q48czpicl3gMvrXweDOy3LbrkDPBW2aPgn0iAQhBlf8RcltHdEnV0
3CnQcK98CNO1bk+iEAvOEhdx0WS84iyjsifMqgaxQ34YLDl30baaxc0gD0LBGedv
eHn+h02ia67SJRgocX8GWd3Ra3e+5sIrgjccNpwJRpVVMF1+PQ/+EOV6RYH5VL9S
+CK/uQyhFvyHPxmZbkQ9MBe2S4q7BAfWbeow35Vhba8VE8pIOaGIFyCsheyWcpd8
SdJmqTRsxePN1Tcy/ZFjj6hBe/l0Xhw0ISZLp+ODDNZnKq0iEdVzn3G8v6VAq0It
ZHRyA5WvYWHQPaQoJ8aUFMPp/eJ98G6wI5z3ePLrH+p/EJD+YX+ffihpSIpEzbg+
wUeqW8bnDL66PXoxKiOfzIiF7QjyjdCyPVIUsB05yQ8VgWM/glKA1bR9MN4eyZOJ
wtE3HFfzD2+W13L6fFQVkwmJ/ErDtZyt2MgTLpcFpxMue/wqfTbVzJ+g9ch+9g1R
8Vl3SZKZDxAHoSCMOo8KgiQJZ+vZ8uWqRaoZLWG4SZt29zbjsIUfskUCjS7/Ghtp
5yKqjX8or4twCBCMm6zbVFlSDUhkXFUzkm9uQiYzI/53doHc6k9M2v26H4wS9JAS
Xis8TLqURfAn5wlge9LGWZTdKz6tO986/DRff0hcRXSPlnBOGl9A55+OEzk7xnwi
AOv5zNJRYGcl4uk3CYm8/NG8/147nfGubUZk5hbm6oUWGDiFRE1eGb8/haxOl+Wt
wbkSfKJVgtmLA4I/vm6eTWFnhRq7Bs8a2Krhz3PEaeOPKl0kUJevBR9ERsPek4hR
6SgFXftS6UIwvITX5W+cE0r0HTUTPx57EJ14Al9rKu1QgqL+B88t9EIkfM6GpZFz
c/hpXCWQ6XSS7QgtQVFM5nQlR0JDHV+UJPdjCzNXcF84jD4nGkTxe2QGfOg54DDF
yG8ZOUGRMrn6LjfVOj+ug7KrnjNbzuiG63XDcIbWg3WFaur+gBcdmrm8RvPQh6EO
hTsIWaNOimu1QLun7/eqO8hacBPKiRJxtspvBxvcXBMiejpRHukpinuDemU2OX0/
9qbnbVrwZn1lwMXIyT4qWwKR5I/qsIGBU7iiUqtUs4An6Y6FFyoxFs6QNpCRNNhO
oHPj9UXAWE0t5c98sntJIdi2h46P1vR8GK0Y8IJerwN7gZbG35o8zmmL5X/KpcFp
9R7f3uRtb7LEt5RTn3R4uhejiKCJM3CmPZneT39sE2Nj94KRQqGORACOzf2xmYWr
GfumRtB3mx43m5biu0kSGGcUX0i2QyNosyNa9dQb+zwsiDMeg8F94CqkLzumC0wY
YdPy30Vxm84/ByxP7rXKey9Qr47NI2iRRRuqvGqaLi1ZmWvznfXB03f22YPEkYd6
eoZIcnwbcWqiRKmppakFjXHvkhCNNJPK9Xd1IPCOhI4ZxCo3bxlr9HjKfIhM9kLx
qV17lEu+3Ux/IIMbAGDKFLDB6vnl2M0Y17K34Q/4UQSCJFOkoUKRIRTFmVLJX88S
LW/215Y+1jqKKOLC2KgJnA7vsIxFEUA24qAei2AbXAWgeevWAj0nD7QUiGbIywhn
j9hMjK81T0goP9caHoFICxzoQDJG+VUDsnPWNVBp6wI0lSb17BGVXPLNeEKXZMJs
Y/MkRvPA7VJpgaXjl/m9IETpYajo/CL1dWjZJ1Otp/x+L5OSknudY3k6z2ywVYVX
dfEwA/bPKgUHNQ8LjiGPckmvnRK0zwdYk2P510oQxDYY12lIjLn1veQXqfj8hAkL
r0wFCWcb7UXkMNmI9tpjg7HiEpu5yCKXHjmh0pQLO8866TwyZ9vEgWA/avaPTGc6
JH5afi1Cn2vKN7s9UWZ8f1yDMIEdZwFG4xS8pYhOKLPvnXtPk7Kicp9qxM7kX4r0
oJRrRpemdP0teg5yEuKYXtne/G5m+pjPIGuMp9US7GRdRGTifNYQpP3JGWCmoUQk
DtktsD/DOe88hGMIXD+k+GgO+By1hPktCBFLwqfe6eF3CJccAi/8hxHoiAOoOz4U
njUJdLEb2FxgsaXOvJIj+fhIqEIx2/9nF+HnC5BmsOW9+rNL4vXI9oGy11zifDJ/
uvupLzq+GOCOhsx98APFSoxNjy6SBiIJ24xSOrNojSuU8XX0UOJcg5r1E/jcKb3v
Oyk5cH6505qxEbgwoObTLS5yMhozdWDTv7QI6jGe0D6bVbqiXsZD22TvrlTqUjKL
2o4Mf7foOmuWv+wZoMLxoyFpA3qTS70MS9j07WFiXlnZ1d473BHzQqf55JL6CAAz
+nUsXQ+YkszlEEAbGM3v7T20q9SO9GtJMqaV4pZ+kZyW0bwPQARD4fvdX2ElwFIr
MUtiGAwm73x8kxn6BiVp0k+1X1lK3rci0Y4nITISgXx/DLKIZqWFKTt5aegrbJd7
6w3+pEQjLXUa2J6Mp8P5wM259UCJCjgD4cYeXX/oh4PoCQNB6CeF8gIoaJvJPm/e
VNKabcnSMiayOFAofe6RDwa3Y9kRKMNJxPc/7P8C3JhPuTjmVTVbZ5Q9dpiy3FuO
PBXl0TJY5EjDmkGk1AEWq54UikWOI2cQWBSLU7MkQZMxvPckt3+AvBpzsBatAhs9
UbOFycquyEb2+5RqiFSCPttsEGDRlkQVmYsqh23w8FNLGCkKzriOXQqfGRifiV4V
Ufqp1hF9GaKCJ4WecD/nj3yEFgPpKbXGeSkz2enKLRIisccMhFl619ePSzcbuJep
NUMznXa0IykQyjC9Hvum+Ff1rPZrcWkItKmAgxqTep2BQrch3LiP7wABxYbpvP03
bYDMdcykCbZg2MgfmLF0WcMi5pr7Nxc23RDINoxdpiZCmFEk7nnVwDxpjxwc/wAy
Sdz04wwKX4d5VMloJTI5GiI4Y+HPbWD+deFXLliiKUHAQMiVFXPlr0SqJb2F0R54
XUqsyp2OAj1jZ1mPbZBfkp94pbwLp6pXyslzGDOqJG47n4VOau0AI8F1ndDWbTz5
NmH0nD3mU2p5OK2ITwQGQspVvMa+k5l0LPJX+A3uHG7KgjxiSGsnXbosBHgpvBvk
CxRlIlq6J/VVyRqpXs/fx6TqHS45YPeSLojkj8DIiIlhRXBvYnuzpnXKWagMVWFp
cTmXxQvz9yJHOnYTEQ5IEfk57UaYJPiegIa0sri3nB1vhEUqN3T9RxrRMgYL00kY
RX9tVEJb9NsIY3kI6AaI2wZDIA7xuujDaSQQpYPYIijDTgn1mt239MV9+mcxmwCB
aXGzmnaPT8uLt7Ojg8tE/ps92dj5UnfBuUbOFRFgMKPOhcRz4eHWDMos9SpCL8i1
1s68bSoFIqeGzUsRCMQJSRR86XoWtm7fRDftYPNBnV3PcRrQzWgMNSa+5ua8pn6h
eumdjQDpWZGcplOifFV5PgwmOIPG/FTq+p6BND6vHFe6CT4pdj4K4ZDKg4Xn8k40
PNo0qJW7ZW888VGP3KNHHYG62vaCBYLJd39bWaPKFnrhGtSjRq+Bk0GcFdQ511P8
jrIIQrTrJNJTt0nSSuXWGpI60CuNdYN9IGDeST1GrgtSLc5R9B860LLfRV02YyoQ
St4N1jX/qbBECidHG4rvj9hpZYOfWH5XUTmZYyOby0XD0pan3Mr+/uEW1BAdrACA
EuIKFCWf3nfSOWs00ROQkZVSH1oGaMWZ11o3LXrgKJg4WQxNki3qxqYhyvXtbi29
fRRDiIa0cagM5W4/zSEEyvussx8ThKTDVM87ZHOLoVT2YjVX1nKpCJpR5+OfFcf5
aywQtkOPoXiu/lZPFq5gqTvf48hLCKYvbSVGb7xqZkKpVL/V7R+dr4VfRu5Vr12H
7sF6gELaa/eKH0rZoSGv7bMDbCWT4rOPKKJui0P2B0/Z30J6IgplSKbKPcC9MeOU
BhVZKp8hRSncj6GLF6jqGVR75xmtM15QlfbW3WWmAl8S2nfa4GG9icWiY6rWqWHt
/WnboJMXJigk5/m797gDpD3eS3hhdSSsv5M6fC0q+Vl70COgxqqqX7i/VgRbu0cj
10yCHM5+xU6oqLnFMWu2+Okm7zYbi8E7E1zH+fQvBPPCWKV5yrTDlN3N6uGLxhlo
UlH6ehGJj0OV71Ab1bdaL98vgAWN0NwwYlObru36i8QDFp+udplHB/KXU57jgsfq
oJLJivM905+rpSY9tR5X4GjDz6A/yuqN6SUIed6vy/efkzp6QfBMcVwbZHITBspT
podpY4nVyN7JLrsRT3PiNmaBRoEUz7Wpz/OA527O2zHGUaQBQbQR5f1FL7nR1iY+
lcy7bb+pPd9mkDEXEryLSjPCZw8kCwGnkGDsMes7hLxhhezh6ww66KGDYpdCEox5
ly0/iNIR8/I74QQ19MAiFHr+GC+hhdKsWk6q9YZHpfF8+dgOmUysUHDrZiNq11oG
9cX/uwsvWrar4CdyNdWfBnr1c/0MtI5PETxLB7+HwE5+GSuYjlP/G3M1jATGHQ9A
p9Qt7bmGvS55bIllM0JM+pnoQUym+NVRL+Pewoh+wYstsTHjPFEg9+Ye3o3E2xkh
TwmdUBJ9nEM/U+rZWPlQHSZhppRgf/dLAYg9/xjfL7Hxu6uOx6VAP6Qb7xOm1gRX
jVHe+IJGOrnp4hPRU0GEOC4CNE6te19n2hOckkccZb1a99/3HF+WxH3WAHbOfvs9
vIbwyE//Y/LjjaEumqcJOLiEiGhuVGSyrZ2iX7ylfAL3mwX2KvjNwCQes2CprJiq
6unj2i2Dv1gV0ZHvcQdi60pQS7ZHCb4iSXeqZBCG3VdQfNcKU6FaGANTwu0kweye
hqNdWqarEXCl22lGjnfeyrZeSF+YMevfKAkyZJGxsKVh2U6AGInxEmpD2nRPm7Fw
nZfKEVFtrbqvmFN76lBUlr1dwy8OrqHyIz+bIovC+3kvRNf7h7zlhhxBEvBv2gpp
ftczmlhDUwYDLlvfupZXxqx2kYqH6kjE1mUt7/b1hmfslRshc44OJH5uv9v2Zm5f
e5X+4Zp+G2h3feeyNUVzMnAxUHw5vKnzRvFbcG9nnechdqdJmP1sbGvk7UQyKo0P
dftPb/wlSXeUYCVrje8zfDVMzhI6xVrO2bf0Mmaxo/+torRBXvxzszqPjNL7hB4i
49oI8aHWB469HqfnV3rlZD2bWpv0aif278iixXORXLr/2nkwfZ5Kbg0z5WBgEqiY
mbCdRyF/qyfznBHjK4De34gCEBprxbYMv/oc3CZtVscrogVw5MGQ4u8DK9h58ohG
iH75c1myC3bQam2ODikSlr1PWVvwTyvPZvDis8EmbUCKgprVwLkuoLzUhkVLeZjQ
BkeO6jPP9qq7IOJ2LO9IJ6FO8hrGGsh154B8IDUOGs5nGBxfR0S/Ocpbprmug/sB
ljFw2IudQmlG1MSD0alhC2JSX/s4fokakFG5VXQi5bDPuHgE6Hl7e2brzjq3b6tj
ampmuh26kXQFNKyZ6YwH1GaPU+vhOUQmvb2bGllqCKKlUkdfUFnEkgW0a4RlIwAF
Fg7tAEpf1gtVchJdDpu9HVoF6rPocxgOVR7lf9KA6rBwHL/qaLs9QvxIDsfioBZm
3g99Bdqp9yZz3L33Jlv+fF+B+BckIirrdjRF0RUrqQlg0cuVxZNAFM8bDELzILfD
+B7K9h7qWvTu3MLvLkHTN8c/RCp4s/ZCD+vtD3Q20o4+gcANwNJax09FaE2ajed5
3Pze87bqn747pasev6btoDAxE3qPEGYQZ8r2f6ZIgnGWVg7Y0b5b6PLbWyEP7tWR
zpRzjiNYLRgfOeQSrOOyM4DXMyFHVO8k1RpGTgwUxtIvIxGKD1nhTg+5Qs+RvtTM
COUHjcYrM1l6WOtqq9iH+ry6K6iF6rWRZf0cZQ8aBLypbfJFgd48GLfuXUgxcoYg
c6eWitnWwTc054yW/Z1vn+eEpMh1pgCjCcTjJGdWgk8UYQdparrSGTYbM49aZyaw
oQxPzjI/anaXDsLUb488DUA5h7/OA9EprzXfWs60V7isQIakTCPuV5YsiPRyi2Se
q0c/uGSPY8owzjwF0Hglpe4dbdXEt5TLuVuPe1r4KGWhqkT8pkN5KJvb1MFp0df7
WtB4P+INpP1bnjNGIDI5T+mEctK75Mj+4P7M4YurFOvzVMwQDStj20ch1GDFxkIH
jEBQfjXK1m/6PUR9LAf1h4Kzr5ksGfxuGOAuqZId7SuaauGYk/LAiAMn8wAQOrlj
+ahT5Sx/sDlRJ9BftVZdAPXFfITbuEpg51aWabrmIEOVMnpZGDYXKWPSmo9ijY1V
VsmPopi+C5PPHbbQnlN2NtYT1TvhEn4CRwX0avjayqhwFYFnnB81c3lQc5IMpdhK
BINdxj3dtm+Puop5y0J+OBAuC3IHncArYn26nMXjI0yG6O5EyM/9Hpew3+8BawiL
qs8C4iVI2bsTgH6gcD4OJosEK7N5VVcHGEBTnaWblhPCtpnwyLC11RKvEvPK2frx
LuhD6/hLitfBcVGdfyToMGn5IiqPyxRTwDMjnt3ZvsoKGkQi7pSup9feKwSSaftX
gn99RSWCshWs0hjrfzfizJFn2UkZ4q2zNUsLs+6FhTWoEPV6FhxEvFfpYEgtpEdu
jIi2YDG1BRMP7pEOUvYLl9zsX5x2w3wsqvOxRt/HvM25XG6wr+hqwUwrUGC7gdac
0dOjQYIweORyY5D2ZAHn+RlcI6HnhNqGNxwqPkLuOlrnNwT+A+aHAPhhsR4PPhft
1Trfa7JroewDpnNxGCkXtjTZy948PjwsFgWpAI3KDPGYmmqVS3XUZD6NuDWeW1ev
nTA0fdTps5o/oMzHXIFyj/oXE+mLJl1F8Y6RiBURryM4Qs3BaiQsrTAhnRN5QACS
+QZft8iAC6YFovVORu4+0D2ylSbaZHjyNNWgeWPuK4rzX9bQ95ehg+FS86KBXuni
vh9jt3VXzc5g32IsO1ZkUD4bS9tgz83zqUprYE9jjSoa9eN/NCeLpo03T2wNZdTO
pCwAs4dpkW95Sm4KQZT8TD3Qzj2KGpRlkVZaG2w8xMQZm6XNL8q8J4rn4vcLGhqF
JWCAME0vV3hZ4oIOR5DGUqlZs1tcODi/+KHGQVKhlm8ZCuziQoeMHxXibPZpwg9G
6LQ1siz67dsylyyyczmlE+My+Zk4Q2Vwpq4w3g6XobTVLUB3TFYsnRXWPmcEbrqe
m4jYlWt0/Oj5hs5xaFDqgAYlaWcScZC/lW8QrDZuPFoK/9Pvqm9w436GIYImKQ24
e2qnKuh04Be4Beo3/SN7Btq95p8eRS0YZdhB9NAyS1aVAfL2Vtj4gDjUYoOrtsqY
KO8gGNxr0a2opdYTtxu22LZ1es9ZS3+D/6W+vwad8e8a2LYBaMuEKpE475CIPlwr
fyRXW7M7ZjGX4tQGt+Cd+m5piJTAzXNU1JJThoo2LbhGpWtZXeUFw05c42e0JR4j
72tGSOJcVadiFowzB/IbZrKmlaSIvFJxXextswWlaFXwepYTgRioezAW599zzOQY
beSK8UiXT0XaJPw/weo6LOMxmANsYbPgk+QZwog90YlVGk4cMJCYxAce0qwS7vRN
BVOkZSTAAIX6/eqEMmNtzBWY5MRHxs7sLgZ/fk+tniOd0b5J620G6kKQVky5Hstn
D9yfbUeZCQSZICr4Lk1Txgtl8m7otoIROtCtGHj33+VXfRaLuYNcgBFC3fIk0cGL
WP95xXa0vy/U9ByRKzIqKO2WtvO0cRi5SvxpV3kwq8pbtngCrdplziXDiDZVP699
2P0taC2CPfkcNKk45oJgaHSWQi1uVvSwC3PywD5VSZW5rEKFdJUpgdkYfFx+m9KY
Jv/JJzJzIxRZLPaBgNro4Cp17TSydnMrIN+8/U3VgIh/GGIY/Rb//MBbj0bmXSwF
JCTmCunh9zO70PuCquIgQaBgZW6SMC/A2sus7fvhartcay1op3qYePYaZ6dq4N4E
67hYtguOojQL6tSravd5H0VjdwFJmBvO5A/s4Va3wxmL3t27XI0y6Rr2KJ0DxQbr
P3POxzikhTeJQUMWKM3vmVo40Rwv9b+5MJ/6dXZEFJGhBpIFmW0oxFnnf+asuoUH
yVXQsMPRDha+WXmfjkhjllKA/z0GYO2iM4I5sOavYW0Nl87pa6qHEfFrYRyVkRFB
nQgz7jPobsGriEgGNvWxefZYirIpb7nETqxab6zI7nALVnUAyLNfEE0GvlyWlnms
DH6YBUPXiAEE1tUvjnjf0fHRx+C/tnw++PlG1Mw+t7TS7HfMj5ymH4Ok6IpHKQsS
6+1zsgNODaX2vGddBjqSU+uZhXIBGHpzrypoUMLTr/YF5cdExGq4FzuE3lbedmHO
E+cvnBGYcVdDsOMB8cGvWAw8ME4H4VbqNihE0dzdv/4QeLRbYFwd4pHEBvENpZIj
mFLwYqKXFCXOm5w2fZHc4SVD5v7qUAqcQgUac6xxTChX1+gylqrDd/IE1vRqIcc1
Ds2v77eXPl/IFg9L+USzgMm4RpW8++PAEnZ5Zs2rFTbk7Sq1g0nN9rRanwXtXCzY
aKDy7QSG/USfRlAXWuYcNJ+APWRWBBjhuovIiFJLsJUKx61wH7LkxEY4J2OaZyek
AaWcKf3tPIccya61OWR0gICWyMQdUcWU0XJ163VU99gy2aX7Y7YtI3NsFR8PBFEM
+g8mQxRYjOB+3oPLEcI2+ozT9QZA5re2JYLHr/sY7jlr2GsHyCqgWtOglgQ4rIa7
5egye1078CikLu2NovK6XmAMo8iENABDOrxLtS78SAtsklUtuOcI1i01jWG8MmKY
WjE2IuQiU9+eaOR6D1JPLKOgE5tNqP3Qfax3ITfqC8KoGUPmleW4kKLqlrQpkR+D
lHJtkxVst0ZlfzOs1RGbjXdBOwSJoKka3HpJQWvlZwUfUi8rkEKPDh32EWDJKCeL
5Rk1acQHQkYhTxkJAveeWi0Nc3A+bDnGpl+r9pRBmYYhmJ6slxoYAwPciwnCSbu2
PgZMQz/ZzkLjZh6dAGZsp+20lodPHL26SdAOhHIHgqzuQ0Rtqut8KF/fB+SaxGGc
OAWHlxlH0DovX2MtzkN2cA9m4nn6zBDHGULxDNdelj8wqLc7zYedzxg9hyPTJU0C
vVvIVutw9kJNlOAvulMPR/X21t+40DK8dXScRLtCm7YBJjhG+5/kDWHOdsk5mgGE
jYgppgBzkVC0Ko6X0AAWkF7KLCt2+/AoPnZ17eDYEF2rpDWsFTtEOjfH2NDvMaFJ
KtKqFA29O71Uy0Bho2brszTtpdn3+0C3uHonHkPQxxwRkRmjBc1YVaNeqNxbuHhW
OvKXTpIYYS6xUJ61obtNW3queYbgVv7G/7To/g5+uQBWoPp2AsCA3bqi5o8QBRBi
sCFtBmfTzsC9Tls53KpndL4Q/83AQG7EGPRSeS/6n3TglsV20WdbtBW3GSuEoWCm
V+G11njEPOtE0SXXVDztrJr4EaFusZO49ObpBTI22c+Pns0KiTRH7vVgMnkiGSje
8pvpAJMUR7vXZn2iN8HWvluj1vnrrJf+ULjo0RRMMtwAL3iSFunQJVcROR9wfWBQ
Tlxvj74l5rY/N3myCfXKz6N5WjhIHtAyX33JwdPpYb10gcbB62ooK4QUjRTzvhW/
yGlehVs5pXTnlTd2Us9HqPypQGfxHOanOkKTG1q0iaYihJu0ItedW8Rd2hBGJh8o
1G6R6E9HBGvfO+r4Q4Mqj2NVuZJEhLmfN664vUXwlxiBNIykMPvWIIQ08TRCT0nP
9pef3Mp1sCe6NyQ3RlYAFA8qL2fRzLt/3Rj8MOYdCl0eK7dpzqBEWcny6usRCFBc
xMda5WBpvlPKO+1mf+4zDExD5e8f/IQV+XlUsh0k+Tkb0mEcmxuqzjwpT/2rBxd+
ZUkme7BOZeEP+Ir5xq5s928XnenqmJkJsJneFflk0B3L7E4NNL4BS+L8gA05Wh+E
jc24MJZ5TKvPxfM+dK7SVwciKoC5QP5WMav8bUxr2Zr7IvHG8En8jDMn+HTlW9fK
bFgo1joM6WzCSmyxfgP/MXgKCrwGgfnC0ICyfxKCgjydKVyShxxAa+MR2yl+rYD9
AYIlVlrJqEf0rCsdHgjFHakQk1prSHntuereY+gpWcy35e3X/w5PiNbH3XgWMI0D
HB1N4pkdE1A1b61cKL90G9N562I2P7PYga+vadSssv6BB/4i4HHrcdsuK8cMEUHd
HJ/hT3plb/dVZpHa1zrZJ/qHA9ruRW9OvdWBKCZ62RPY+UeRBu5C618gnmLk5KFq
3buLtlIgMmkJMan1oP1ottM52VOEKhPQgvKD9gR6KYUNhIDdA1GVbFZn4od3TnHB
PhapSvr7HYXh4m2nKQ692c6iOwSieN+1JyhWwVuINLBMjQ8yvaNoWqmnLcuz+Yaz
tAO2mbQDIlcpXRVXIWsA0EVe3I+aajyVXuOxTSMONrwYNfxKhquC4BZfmUXKg2KX
TXF9Igve3DIP8T87594hDml9y5WhuJdroktuqTaarBxl3XoymS7MOf/roIqXfYHS
4V4njRtwag0ZTKlmEOEkt4W9yNUrv/jEPLulYuHKBQ9bXa1B2eNv25MbWO8l+8k9
j2+bdO4SEvRUDaOHTWcU1eFz1fYT4m7WFb12l6e4U9Gvo4+GRrdoG6TkeaqCDiOo
coo/CSkh8h3KTeo3X476vQKdEL+ZmwqSFougC7FHahJvGOJNcPz65/SY5+XLv7pd
mZmQyiuiEcaK63lLDIWYWMdoZKnQxWl2NPdkFXJtJm5HshHW+Asd03zAGnJz+Im4
YwpGcw4mQOBXhdEaeWeo8bDquWvqIc6xF0/7+op2o/8Hr2p1po3vJ7Oa2IJDktOo
+sKB/t7vMc+wlqEp+sVwIpbz6MEcRfTVEGgNIFTnNVoLHR0cuMa7CMaEa2u8X0K9
weN+yjeq4p0pA7wSF8sNTQdxL0rfMxfLorn39fsJmPooFq1zcpPHNv0uifEiLl8v
7co3K3edRnph1cjIFJJEU3o8egyWxICM6KQUHBTMrmjQUnqWf1eRwpu9Pp2z1FcS
vKCDJpLimUzxhcLxyPJOWqBR7DjG44Rmf/8Tdx+OkNP/Z6ys3v6ZcongO37TKfIj
dJUtLeMB4gucyI6uxx2mPIZTleVeNglMbWsuXmzsAKHjNcwOfjVqopRw3ET/Z3aH
WIvLwHM4rfPNhgtAIOKXYrxdp0ybxAB2yF0twMv0IJ7g/hjrs8scMiJReRnV9pNQ
hPpZOEJSA3mY4rf1huzxiY9GoagfJxl6T/WRcY6SBYStQfUO1FtCzypgMuNusako
pv4S1OQAQTByk7jA9V0cG1CAO3NXAtY5Dxm2nN0e5BaRCnJplMDDf/orqKeT39ce
K2u7B1OSSDmY3DjIHpsCBbJ5klHGWCO8edXufsPcc14RMLsQhxAabnPRuz9O5Pgb
5o5gAU8UQ8HWgwGlpRcD0iS/RnR+ZdtMD4arz5x4J/MoY/y3GjZ2IiGSSM5tAWSi
fYHA5u7Y30o5J6S8GZhG43U4ZH/zx371p+XBCrFaK6yaK566NyC6Amn9sCMkNaUw
67h2yZr9hitbtR6tdRxrzkVrp3wwjGnpQSdYmfNzNTgRL4a8FmKMT40w8inBHOnf
yiURjoWsKlKWqAxZkXorOf5pLUnqP0uL9d6CEvUCmYuF3RazJOS2JJQevaFMDuKx
87Hj0/xPzWNT8fr8KDsbC+5jSwEpIHAIo1UaONZMF8/ozCcJHabc59MJB5Ye3moB
h/LD2PMoHZETIjBmIQnd/n3vbdJ8VsCsLpnHvGX70JzLuUN/e42EkVwZINhyZmz+
Mkpo4xMaq7q+6BqF3YfV7rDLB8IWc0P7xJGmcR5gr+bXHv6EiqYaRaKRJgtsRI83
S7LZhtS+7KfUU1TYTA8QxRLy0+XsXBeI5JzLajUl7gxDJ5UX3zqWzv3Vej8JG5aN
dhWltvZqKLamZXVoQQk4gHVeah3K67DnzATBcOsfqSEF0qFMbnnyvZa1qPze5VyC
f/1jrLTolpVxrr2/xbptjABtfDl4DR8Fnavz9MXoSBP9PeeLUtj6BRI/YD0KkYrM
lSEj77ZODuuP6yCIHUCtm6p2Nj0to8Mb39018NAElJWa5V2Nqc5Tg7FOxYSID/pq
VSm+L+k/lpb12JgekZj9uU6hEzCuc4/8CaFKyq4gpzyGYuqR2WKIbj0szYA+vX/G
nQC05i7VJtf9sDYw34OaE9rg1tBfVQAQhSZGIs0fkFqEICtZQBv6bTqNEjzh4IF0
9AqJC3gYxil01dohU2khR1W46bjsN7TbTwEwNJjQd7zsIR0fhDkdaTQQsCnEwl9B
TS3jdmmHiFZXKSGXNb1nGmD7HckbACIIZdUfPKv7/h/GmGX8LYr9HqBJJfgKBQKf
Fw033Cn6R/9YFq2ElGbdF3I2zhcmr8ebz9vHeD30/Wuqx82rro7hvu3ZkyJMRANQ
v/Vzog6wmpp6DCj37M31qCpU+C+nU44zRs1p6lP+CmGMgRPKOPufNvBAe0yMmjnF
WSYXOa8hyVUDCAGj0f4sRaQfis/0nyIv79q8vf90Lcwe/aTs2HUHZj14F7iUrndW
RmimlJgLo/TGyYnCqu2iWNCvdfUG9Y7kK2EU9PRsZJN/w229zKc3OyyJVTL5ha9E
+kazTAZTm4PEzglizlif9qhBCr0O5L8MaKz5/B3wE23FI/2d2ypkVlrg4GZpR2r6
6RVacDPMg9nkT+UXrd4LN7nLeHLCwbzBLVT/FHJ7lSXIz7Y5UQMeakO40WIbyJg/
0CB4HR1ajFU6UITl2jj3v5emrcMrh8IibBAfousrs3EMZJ3WRwoaxID45ldgqpBd
O3f/W04pUO0Skl8tI9jZkh7nSTRa4ONXESDXovkofJLmkm9C3PPil+tuL0uvDJ8i
yvQc1X7xoNAiTWqUzGPACnvvxz7WplYdJ4ixBcit9fiwtFI806kDKAkN2VPBIQKV
/qNWiI0jJganV06leX5uOW7Oh6TIeUuN4QD587RosaSvMiW45rpsvuRIlBBzwv+U
uzbyjZ17NSDTP1ycGjCEogyvWp6eUFpSVR8jv+a8NxfxcvW4WmEik4Tg1wPfakW5
CbFphXk+n66SrnQQRXLiptlSB0uPkf5KLYpZZ5eaV70ujW7iloWPk5hxIC940nbG
aP5P5fooCuBqxuX8dwCg4HyqwEkxBzZ6wZDQGUBnINQ3lPP9KD9b4U7mNUKZx7Ri
lU5tL4BzBShb7CFVgP7EwQxlML3THBlnI4ryYrr46Zd96Ax6YPCztkic1P0Akc15
VfGJkCI2dyvMzhWYTmYoyQdr1RbSIxjuQxuSa43t9IBLzKG8OH9OONDglSvQXI1L
ElFu8QfKj5/EZfwmjPg9an28H0sfZnfBlqna9YQFvq0dRCxwCSZWkcnvYGZ2Qp32
igLtH2yS6n83nevYzyGAKnBMZj0KJFNRE6VuVR6+WnkkYM8uYG8xuo2PRVSuUthR
hil5c99/6jIe5JcBvFAVY6VwyOu/4jNr4n2Eu1h3XVwqfltXbJaQ0AWvuC8miwjT
/KbPZQ9jRXyCkN4pDEjjCVSt4ngJQG6phNTmCWzOygIeBEsfiKhmxONZDTdOF+zf
a7O8PaPyXYAlHMEvYryv3F1cl/kj5sWO8Z40ay/7MbI32BhZHI5PZJCI0snlIX4h
jz/wuDbdhu8ln6e3HbqAL2VkKv3py/Dgf3Fg40kloaLBMvmsVNCAinRYKbZVuAq4
DgjunocSNPESmCvgUF++uCKYCwsQZdNkmvXeW3xCvkuPXj4qYRQ2JH46jVMchMF8
19foCqApdKp1nZ8Nigijz1aS0/h6HEGC99DA+EbbM7nThTsu5wgOZjhWCvA96Gfe
uMYMelqUJfz+69CD8whphuYqOxFbXEghEp+K1ylV5QQAs7ZMlaY6zsqpCRcSqAmD
kMKo/aDqZEWH33zAzAG1MsbmOEbRcUhB32kkMrGhYYRGRUnuFg4pxX8yc2lg6pgN
xO+PnGlPmWagvS0qeyhkhXJvSFe14hqPbvCt9dI2S8QWwpE4PDdMeLR6l0jfoLSS
KgF7NmKhsBZTVWSCYvVRU7LjptcgYqxJ8BUNg8bfDKQqR7VWokTufEG3u3pGPu0V
Z7fWykKVcHQ4pY5iQTwzbti1tqIXMTtcaMOmdDD90ZxAhZt6ZYLRBJoMi0iJb3sW
HRpHXAZjcZ+6o1E2aSYJJGlzce8aoBC1yewzPh5b1HKQtruBmFJXCXTvdzaBcXK7
B8BMM0Y7PkIaB2rc4GNiCqg1hmKbsgqwlP/GklOMsfO3fhnvSst/tMHbDrSB3rHu
EBJ7kjxvG/OYMgTbx1RVqWGkLc1gv8wbwos/ry+85M2mC3i+qOTDT+D8dohYs961
BBaEMneWipqJcPMlIumyXxXmybHwiviNZ8QsqsR9q6QyeL4rouQBogcndn5425iH
Ax/5SEVW+NXn6AiNdPelcGkV+pgfTU91y6WSYDdSAacm8ZstUxwKdKPXgKbu9jd/
oo4b5FTtRnkVxrerOfunqEjgERYkNO+ZbcjYWIjl83kq/sHGWqxY03qst6O3Z8Z+
UhnM+lChgo1q+At36v08r0hkcHbqYtotmFBmtEwzOSjLk1aFWIi0Ug+NKhV8Ad0j
r8hszKC3hNqnBqucNQqyrIrxRvp5txJVf9jPgUjA9xEhqFHlul/Q1k/BkBJ3/Dyk
STQijlogfTiaKj9jtTx7iA1u3XrXv1JxLpOs2Je6Mv5S8l6mYwIHxHZUmPGgemwC
bwhIV0LJe9pSI0E3FudkHj6R9gfvji6h7hg1tX/b/uJu799S6czfm1IAc7+jdGUt
KyZNJypVe4FRuQn+o6oORRIXQY6MCVIt7MDOqQmtZKpl1/WUs5HxjtlDvnKvOo+q
WziqpPh1kbB0c5i4KMDnIe1hELT/s5ybr5doZwjQ/wZKyfvm42Hqqj51VckY6+OV
IRJyQFz2raFMqm2wOA2WMFw8fQMq5Addzp1D3RjlkuBtd3CyIF4rhyvKJI354Vcd
uUIb/fP4y9U8xdN5KsUzvf8iuCAnzhHbkq39p1k0iyqhKPPn3jDO+/fTKUH5wchq
jNy7p1d18f6KloA3vKDoU932fD1rLOc+BEjuPK+0vPQLA4F+JSXF5xhNFeMNw/4e
iOm6iBm7rkurb/xC9euN2eTyhq46c8GmjZ72q6h2GgEVaDwvJfQhxpN2rkvUONUG
Ma+bXlscT0aGFeXuxz+vUdivEW0gMmWAND9ldxMqbqWiKmiXy3GGbiEZ4yo07h77
LwD1XLZpJ2A9AguSM0QaXAEmtQAxSHBGsWlp0v5YaZf82nIkBblMIB+kcQH60Zq5
G+L3oqK5LjnYpVKRRC6RxFqMiCANaK0ICc9zIF+QgT+Mf0foBYPlCNX+g0SaXiRV
kVmGnVB0TKHnTwibNUc3OrqwnZDoPhAtbgpUqC9vQZEF0sxZyJjNbn0GB6/7iKrp
OUT73hq58DFbvkmJcIpDRthOhtfdFhNb1sLusDrX0SbRie02/eMQs4VelvBjlf1k
EBq8kJS5ZrE9C655SvaIZ8oXPiTwCnzfCMDqVlnfJkjSgNlFM2jVybb8O/6YZbj9
mfr+tknsgZE9g4jhq2Q684O+RIV4rXPcvFIu84uTD1DyxR8vovrYKmqIw+mfI23A
BM1Wf84Uhd7juAreqfWQ6iQdWIJFpK0Vq2tLvr8MmZxkypGi6uAHnJ+Rkst3Aqbu
AhAKJxuTPhnK8nuofDEr1e+/xt0P+F9/6qUsOmn9MHJj/sewu9Zjw6HbpjoDmKDX
Eu6zhPYMj2OwvO/i2InRHimHxfmMwhH2gc04AHj/fTGmJFXFNT1fC4Mdm0gF5w+/
ALfsjBhaqTaYmaP751O1yMYYfPbKyfjXkFQwqxqTuHowX8VZczklWe8pOpT0QE11
DOdhZnpPPN1JXF5Q7RnT5O3+kHXDUcjQEjgA5bWqvi6eWD8Ua2HitB3ThTm6S4iI
iG+uql59cUQ7axdmMx89VTM3oyxRLwGdodQmXPHt2YTpDAc0TtDX94j8Z1FXWxbT
dk7QszQjQWcEIWkRwQwBSvGVjI14sl0VoCICJD+EYlRGc25s4FCq7JJmsEBf9wPz
0MJHIG57pZuyZTMqBtjpvmYr1HL/8RJeagEtec0IOJh+SDLAij9JJz0rDh/ZsJKf
oeOXpy2rxa5EJyzi96/qNl9d3bbJm4g+ynRSwYeyBzs/zax7RVoY9uBEAJjbbFSU
rD9ew1Mx/qMR69IxQnrC4hh6q8iBurHDj9wVu+XwV5ZWnYq+Hs1jhys594j0eGO+
rC8s4K6c6GZZ+mQR0Xm08y6K8HJfN9QY23iMob1Zh3z8zMHRMrf3vXMnVRkNt8pW
OsLk9I3QLVD/tUnTizL1yms0KgHbhBCnV522kntx5+YBMU/KweQ+8xVgQLAWcIGq
69xwNWzX2GeFkwO98WUo8UIFaH3z8SXisE7LVmyl/7df9DFjd/FWmnr3hLPBDyaI
lo+N436ViklMGYsVQNakxQqnjZNCaeqp88zPQCI3Q1N3LVMVw6UOErx4SLVudxRQ
EvNBzAJ0f+yf+ijupt9tg2xYKEu3++2mO1LEs9/jBmra62FwGk4Q6wwYTOJGXOk+
2PqEUuW7fSXUsCwlPoQ/r6kDcI9TToG4j3rSj2W+WypLdsKXAp251oOHv85Z4xSj
axI+tiTF9aYcUJ3iBbzovfKyAsTZC2mBu+VEJJHC0i2TB7VO5OUVwJGF8vy62FyP
YGx02bRca+GEweNpSYxxjPi4s/lixfbwYRTV2BTexq819bY23+DxBEoApj6Eodko
1XnREtN54Cq/4PqCmvclSvruJ6oFmaxNUxQR20lHa2zKSCq80XMSawanZd4pPTzs
Z9r+L3OAhi6bQ923+pXDAb7T306rnoLonWHm4GV2M6GNofgfx94K9bqKd9i53iTx
DI7vHV/uWA9YAZk5Q6uDxlI4CdMVeFvxBROAhwP7zneuWVn5SfXF17Eax2fg190o
TdcXZPog1/hdo/mJZOL/5Hp2gF9m2/bgmYGTzdxzHz83cj0I6OBao/wYNpZx2f7q
o3MRH0qvuWPJ9HB+M1Zg/l1S7aGSMU0NusUqMN5Bm2EcjTbi1HtAOPxVtz4mu4bo
uJ+OmdV9ZhbTnXfk3rzB89qElAILYa8Snz7y2CDpXky+Oi4vcAdavboXGIcCseQ/
addQ0Z/g++wYCHjUYfPvev0+I6rYaEuY7D8poJy1q4pbNdw20M1OclFCQg39JAxJ
`protect end_protected