`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 41760 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
S993bpJjwxtMDn0RNN54X+vne+zl01hRRBUB1Frw8nJIYhO43Jkm8+19oznvTPJX
FUGldQu3zWrNk1kns9pasXKnQK5az91G3fGo2GVk3qsGDMcFgPBLFMpV8Fj6q7ij
fEWHQFj0GvnlTEVqVFz7sKgAIa1BJHetjKiO7EQ2nqXdDF4LdG9RMflQeoppKK29
jEaNv6+OgaomiDUSPXFBcdPVps5jyiGp7dZqDl8Kei/WLLD/aA9QyoQhYvqxi5NE
S/Twlr5uh7/hA9O/rAaFmpGjOuPjm2ZQ5H2bupvyQmH126TKza7/2DwUw61V8gBd
4BA8ilGtv0pFr1rphJfZNO8nnN19DUCzBX3xDCvj9MfSaCM1qPermOPFiSiEzkc/
g/Z+yQ2q1UqVIbISdgWQII+inVL80ImmWSu+wENdD/Sbo7GEO7TraVMKhLGUcR2n
GHe/c3ArPjAY+G8d1+zNiALjH0mH5Xxz4n+nhNyV6/Evuryt7AzVhdA78syJHlw8
kQRMyTBq02arut33lqMQeTTrrZeGvIvIbwSBu88VLeQaLLEiPmvA6jA6r4WuEBmb
cUnhcgxSCNnust+sQIAI3003/bJBgcUkv2YTe5mLnetyVAUwBTbeC5N+n9hT/BcF
p1WtDj9GuzkGoqgK+Icz8oOt1ky4gjOAUVU3hTSCKf3djNrYFfVo/5E3CsEl8HSM
U+S/HCCFFwO0xf+U4xIrqOpcs7ByCi/C+MBtsKB9v0CP8jgnJk0jJ86TReFmoN3D
+IoTIXMXT3PoCSRyqxw2k3lYL71N4l0zB9F9j5yxLVcpQs0ykRKNfbUQr87wFl8b
FSvaeIrptO7fvVdOmvDr1sTdQGFgdNvFytHZ/nFht6SWtyl9gy3RigPLyTEU3BJn
os4Y367/j8kbLfNL5zgzqCfspVwkWBHergRzRkVMxvAqw7oWfMKpQps65rEWrCuF
IA5gsXIGvxphcfJvVI52rcJZo+vDgpSUqjpdZEpFO3vc0R8f6LZpW3V9tZZqzkuY
tzukwplLQnQO9jGd89ZBpoOYhytMS4PXbZF62oMGbWDseeG1O84vGaaoGOojQqgO
tKIR93fyOZeqpMIFiWr1x5F/de0ApYKZIRPaToN33NV2SFJZ2w9cvnaxrXm1KwsS
lUyUOm74AIWktsYWAfC8RvjxQiFotRIJmNf8xM4rLY+4BMam0rbTsnglsZcy9K4S
rpC+mi/Qkc5BgBTfm+MarAxDk1+KEK4a0Z/9x7zRRYUBnvff1hBi9E4XFbg9TO2R
qcT3vE4VzSQdgU0kl5jLrtnc2SJQSokWzCG5ygNmRRrhZs/ulrEN3m7RZ1VdE4Cw
pNOqCP+vFg/GC31dQGS9Av4KXYFhe30vtS0iLIAfzMg0yJ3gH4Q13+KaPwgG9Znm
rHzTl9o5fdzDt+6tmG6YTJYH9ao10Dm3tp1vUxYiNe6p3NAFIPPX1XdPlWEP9xHt
ujxRbjPcXXXku/T59btihCrE7AvvA1VV94+D7BMk+lFR8cJ4ZCMOfdblx3I59CZU
A9IF/LVYKU1btcblr1DJq62a7roDH7LaEto05M0nHt3B9z9/oRurnV4skfH3QFZB
8BCuyOid5PjrBPBzXxCF8eOCzNnFvBGzVFVCH05N40KCJCbhGGqZR7aGMwF7LOj1
rqBx0LZiVVRHAUodwA/e7ST7oDnyO59O6iMBn6TNiN4zAzOICZZxe75hv/j9bMYf
6HLMVLcYtuRaY7W1viJyXOiXwSlFD3pacuGEsdTw5JUmm70hmI5k3HTe+Nxklc7A
AG512os0gykZxkVJhX7+oSN0Q9drWczD+QxymGxwXhrQsARZDH4YZ1/qZruC3DA1
vwLDFwW4oqi6asC81zqGH0bUHlV3YtVwiz7lm6UBaMSQSdaqxi+Yndwp8mo3WW7Z
RBzADqRl9gP022jrzOzf9uZS4dQc6FHxUZ4yV6AKGK8vQ5w8ImuTFlsHD9qfZNk/
BHesAn4KX8WXnNOLZPx1gDzspAVPBOTC9gVX+Ngqbtc6qNmtfnkqRSydzf9k6YZk
vre9jik6bpMmnQ1ekf9fHAHIhMdeYu0b+jJmMeAllBZpSWrwGnFv/AbaIPKYO7/v
npVgNF1bbBQ/AS+ngWHNE+3rHq3KJ1f1wPp4v1QzaJuZ1tNx9bF31G7TrgGKPBs4
QnRAa9E7T95K6EFOssv02wVupNV1pKBCJbiHqY2c8GZcdyFIBHtZsveszY988MPO
kymMcu18udM31wuwRa/XUtAC4MPg9V8vCdG3jiie1mJlcjMsPmEq1kfKa4TYAK6e
Wr91neQRV8Zg7jIDS1RSVlSoJXIJdZy9weqNRcyfPzJc1XaM+lIa5A+ZB8BFTnAo
HyH6isxv6GRr/o012qiH+2t/yie54PQ05GRqhQQx4ROZxDKNxTf8ZA7SwPC+zuUf
CXBwGTA5KvDULHWnu/hxONMcrqdTvZiPAqWAgzqjUSq6tbdZFSzbiBAwuPZNs033
iglOEgJeZvPXMaT6U/qfzCDmsJ7Ne3/5xIC//AjO4C3zTCRMG2nzbbkfWqa937oo
AkYV6P5egw5WXc18wm0uNeOznwssEkWJrwa0LPJzuGJf70epPrQU5VdeZg2GPgSt
rlVognbECWP7m51lUP86xWlwfdQJl08U14Ix2EgQMYyq5oKNpZ3mE4e5s5Jg0h00
fZnfJBOo9XkfWCt+k+xzUsFdNzGnCtme+IJ00h/YgD5MnBsR7DOPqJ03WVnUK1rv
ZH9nL328qImh9Vx9x/yqXPQ5/Y0gA3BTN1lTtakKIz2JnvWzjkUZPv0wIcFcZG0C
E5JYY+S3Hwra00rVmUSwx09PSJYwMfkVHv+9Xghm9HFjBom7ImFIYlK46RED6oe5
8Cx9pPHOuI65unDkdGTSU0JkTb+157/XaAqN/0EsfjOZukJcqohwdZ4NQiY+bKLz
p0G28UUNPCi3Z+Y+sg5aFJllSd/k/4Il1HhRKUnHSCf7LdADRcF5T6++VZW7CMoI
7PQRhJLzxaq9kU6pp3fwEqbizFzAvaIYKY/APHVCqKfRVbgSC4QFfLLUOosMkyPb
IvRUBwn5uHfsO/IZ2ea34In9q5YW2hNu4z/aYnyfogKG4hAy8yur47mqf0Jyuayh
ZvbxY6uemBiQtX8YTOOBPLnAezgb4VdoA7Ga2UjpjMFdRuCJ6nMHN3mSlS3u9ODd
SLenIfwToTnI0E28jc/kYoKz8vx7ZvzBTgZhCVI1d6/MLtx/1HVDijPByojIM/9h
lQiphZ5Mh1UqQwt+e6uonc9OsrsFm8m63W/6kQrtyJO+gBRDrjALLUQSNO05f3JS
IE8PFpWmSkP6IHdyKNhoIBDhis3lmoO5kA9mbGrTYIqtzeN8OmryE0yF+m1el2WW
78CdF+HRGUhLF7lkhgVGT7uHXzqVxZNDrhglIW+H1q14ac+t8Wag1Iv5lxqo5tKO
TdACSZlrYIANuQWFK/XlWFuY8F+3FQlOfhUVrHiAneENa5UIi29rUGaKw4mP3ER9
mqFWh+IR2hRWVPld9ABJIvM1n/mI9qZ8K9/orR06SHxT+Ykuu0hIKOm+P+nSnwG/
0g0OWUdzxvItUQTq6IVQDFSwZlU2satHrVF9eWSFQvsZ1rTNVDZbYuYA7SrcaWj0
nf6rOWlkGTRiWf87gdZ3utBmMqkekCRSYs98StzQOKZh6CQKf+yH43iFrlUIA3nZ
ia2OWsJgd7QNSFSpfbHjSKUseYylCdXnEYSudU1Vi+S0yj34Eo0keMP6NrhgETb1
OAMntsiIL5xR7Zqx7l2pEWOzL5KrYlFYVK89JMd/r5m8PMNbOwyX+55ZKZF5ZKRU
KBlMlsOMQ5mjRrqFcPcH37XiyFf4AnGFyWS3wDgpucYnI14tz2ip2MQ85zH4nu2S
JGwcNS607hc98aQj6/wh2Bg92oZ0k4HOTQmfYyMfJqSotdWG30mGSgxvI4m7xFUg
7jK6ZQPu9Cw3w0qYtfsWPgHl0n2F3ZT68BiNaVhVpYVYQ9akoDayk19UtXs9cetO
CxxXHhYIUUuCiPO73zCC6WWY6H8kukkws4D55sr3cLYiqOtVdNMVK28VvRCLdRgd
DMxFuqkFlxGru3zbDjSOIsFn80CWG/wiTbll2//nGvSNvAVBMIzNwlV5fg+YsSIz
dVrJlvoUDvd8hexti0ee6GhgyboMfUmExqpYK/FBRLQd70yW8V4K2LXBWeeaEw26
KaS7c2OfrruKNV+sm/En5f1+FCDf5Sgj9kqHpXMW6CUVDYlIfn8r44kZhFnsO0hh
y+77tWzywADRk1BVLxdWs0jvOPr/WOlqgXe43bd4/R3w8J17jgOUIRHlx+SPziTy
/u0sDQ2AnDX1Z4RADmzGCR52YeSwZ8HnQUtveSS90i2GSaJXgWt9kiiYlGUqf/FA
9aAW6kj1F7WDYHbbBa1WPXHayB3bSGL6tZ3jpbFiyqpXH5YPCCn+RqXFj1Gi8Jfk
zUe9+jIi2k6IpcmYjlGIsVex2MbM+TgVgzAXtO08cUUVu8UuSDQlf+5L4x8txh1F
dea/08eXoq+W8GX4Gth8VCE1Q1HHgW4kqJdvexTZdjprjLf9MZzELW/avMI0NHC7
jV8GIEULNJanxJfXiwhVP/zfg29lLlE87Zd4kXIXTmTKkYD6kVNpBSA2KyNCTdyz
wx2AWz3NvaNPDV0OmXFcRP19l65Tzho/CQTPRsxgn9gu2vUN/g9Fq0S0oGQn73q8
fXzXvSuIbdkcrhTw2TTygn1/hGqMwAPTVKi9C8zCPC8XvpV60pvf5vDk9Lr1YjRz
dhIBkRMTEvXccc10haHpqVDOaBgJsclzSCmqvGCn90MUgSXWwhZYwL5BQgYsWzmz
P9c+wSVdZSbqzX93QtulTzRlCIpTBQcwcb9fGliHu+90KzzVE1oyX0/b7OPC/snI
97DzBQMnfs/bxl7v8i717zG2uxtEuU26OKjP7eM9RL3K6K6v615C9sOdOiGuz3KQ
pf5lcxR1NS/YeiRKnSddvovpWG+Hf0NS5AE3VHa3Qt6PuQdfHjDmGMdE00uHruq6
FH78b/zCBIyCYZ+CPkuhwjOLZZyq9y1Ilrl0ec3UUENLwQq4p7mqNgLwDgy132da
NHsQAYu0j/jn6uwzrgnAhTC+SVX2L/XT/i5JkaZWBP9mb9LlFqEVuBa1YCBndSgJ
XW0Thl7wC7dLhUrpppNfeadcejnLlYW0qWN23uelidnNIde+kdAaW9z47a/HiGR7
nIwZvSkJIhIzE3JtTRtc+gnq1hbY/DC/BQ81AMLm1Fp/RV/JtaAk8f5vBB/VagS5
qWYXhY1asckX6mxDzCMmDgqAIpbSeRvNi4Ljz5IN6LXpuTHCNRmrPCIOo1IZRFmS
XmVg6OHdFw24KozKAaYeq18P3fLHnFBgMTBW8s0t2ynKMeZcHI6mMj/Xm8C5sPD1
320Y4tmAtvq5McmatAryYYp9Gw5MAB7Fvr37pgKgXrfh4VG2IZxLHs47w6Ii8TBG
Tq09IHl0ZlbiFxfFhJP/nAshBs0vp05zTMANnoXSVwDB3DXHtOZnW/IcomxhCver
q2TkKgBN2fe0jGjuLe3MWNZolYqvwQwDUS/2/zpeIUnF71PGv943HtBVzEd2a7b8
kx5ypAFkDwYw7/un+Rk1qQJEXxyFVtGVnQ/O06jVrRqh+I4ac4bsPkN9cdKJzLNw
DitmFV2i8GDKolnI+ehGdHl2UmxNg9WmhwrIUJO2F6Eka8g1oiQuNamxKmPoDEin
Elt3GMoXJ9h7f5i5yxv9M78h8xnnC9MQsSooQPCUWak3NKp2nstsqllbZeodCVTp
pm2Y8nQsxZs1aWcbq5BBShkMqqGOUkkrnXV/z3/y4aBeajJB9fktqZaiWle6xZHf
FaS97VRtSox6K5eWx6yv26K66SikSceF2uwwnmzQbD5KndHPRl6IF0lQ+FryuhGU
aODduPgu/FjHFr2DW9eD4HnS6n9IQ4N/fV2b5Em47xgxuHH1Y6exmrLbfQY8TliN
sI0YjWlT8ij3ZszKFuw7DRMWnqrTAumtjz4y+p4RPhJLwHrp9h0jXODkRq8vEx9a
rAXS4I8OiGmghoDIinbLuK5Xxh0dsjT7mev6bj3QDsaOQihVz+zwlOykqRQaxmFi
5UW/mfkXP2PdoDKWx+dRIxFPbhjsIrLf71umFNP+Nk6FJPWkZJFz4RYLQtM0y7uM
3tzBw6sUXh9VCICksTW8d1S36dzJ9PL+I01hgLjBwaAZqg9BWu1fh4IL+J292LSa
LdOjTxBiRJZUeELnoV2HvYgXbjK78zC2jiOG3tXABinERjQ9u8MCiqcD8+5Jg7qQ
JXIaYGgOaKt2YPlGMIGWVN/EqnQYp8MI8GK052JjjlRTt6AjI94lr690if6cWLj9
Uh9WDjQ9hqEBkmdtk4ma1jREZ66Cebq9Jl/U+4JaMwU0pkVxDU7rVbvkKE4a++/L
nByQj5Yo5BHy4sdbxevLtMO9+xMgXLWIclxXuoygNdAlVa3gjwbWDBy0KXVavoGk
fT6g/8IP8DxIgXCcDdU8ykqRFzll2CoJC86ST/NHPR7fYacYDjxDOl2I4tJe3Y5x
eCy272HTALbuiLyDWyBl+71l8sfW+6JaW+32gyD9/JF9oEalCKipeBlKC77G9bvR
SSF6jgmWcoOcvziR2VRMYmsGkOUZGdHtSFBrQredLoG1X7MLFtJJINAhoGjVJ1z6
e7bqZEVGq2Jnq9q4QIOULiZpGtVd/bZidLviE4lrbr37U7PHvLJlMT/89MwszpXQ
RpXXPiG0xYX/3aDR71ON1zaVbdQlmIluC04JAJ5WaqhEpKux+VXrl417p75p43Us
fmhgdcqt8VUNDIo3NtxTVJEa94b3TWnNjIOzi7SrnQ+H3A+6xwvx9drtblxXHPYw
hoNeIwvmSVNWtL7rgbRzy7lo+ORlpHc+3YXcF34S/HJ2LHdlU+fcONNnRGsyB7zo
QJ1mFdBrYq13gugHZYtgEkIEiWygbq+/jNmhrrAt7M1fUpZNNGs9K5zF6F3DMQYO
PEBo6NK+EG5s0xOkZO7GfEzlvqukXEG5kqQ/hOMMT9c0dm98CutzBO1jXRUMLsh/
JGwAn2LRoVgD7ubM01ECAXzEvlUn2NMe6ESG7aT4+VFA08zHvquxg9Sk01iLlblj
MAwGrnJdCI4+920i2noMeY2ls9okbB3qR6KnxooFJdCF4kXPueWRPg2+AI7QILnY
Z6trsNcAwSEtSb3rnzlVwpOQ2bvdDCKDQlgBiMDRB84I3RLgnrqBruHlsdpDXlb4
IPUzC2XOvdKzvB+R9/H8jZE/EiN/GYwudyyx2I7TVBhWpdgjSGqm30waICoJhzmI
1ImDIvsGEDiADVp2SqKgPbaVDqi700a7kZHkg6ysXngWf6wFjy3dvUVM7jBkT9vI
WKCjB7N6NXs4MEpXahesCEn1dU2VJ3htlDt4JddcU3/jBxoQ4Up0Ba8sP56H5s6/
IX2XcaB43Sme9AM/Z+cVYYUSQ7sUD1adJTLi4bIN0iuVYkA4BrWZBHp6WSLMgI8w
nbaqcrazf2Mgmb+QHOQWsij0CpuLWrXIuV8f+nJgNvva25zf7DQOKGBZ0YBbOt38
ogWoBgKFOiUgobBU1O1+8DUiovdgdMQnh9DS3RAQm1GJBHjZtix61HEcA05g3b9P
J3eGkT+oKn62c4+NbuqPvEw3viUiSkCyePwuDnIQsS+CCV3AVvYlR6M/Mc87MGbP
mAI2Om2f5YyjuOX1rc0hqsiODQ4f+YrvHFWtkpmWCYYbFZiw3xTCG8XiUdhTckAF
y/4x4PEWAcNyJG28KGQH/GolUUcjvFq6JgC5XhWWG9E+ifVfXBo+WL3Mp1VU9xun
O6wLC9fFUM3q689TterAk8cVPsscrkBhpL9W+lZQJG6K+aoMlLy7X7xOGyhKtpAY
XTyQL34f12fN7sYBfPc9Xcq5nwjeIpfJeN9B81Y0MhhhM28U2tDEymbxLqR01K9/
4H6r2EqUDqk4c6oN39z6UPvpOTB/1xVPHFF9+GwRy/A2bbakSoc1Fli6JYQY12dF
p+QE140Qu1yX3CfgSZOV9MV6vYpPXFkJGlpCq5bviHTcYJhp2omjUC40tAlR2R+s
JXYpwl3AfO13Pz4lZIDes8iwvRhV4poE4W1BOWPwBN8T+mxLUKpvO+OyxAhS1bRu
V4e1mHgpZGD5/jnSoXDfXxbZvrfGPKaqHM94UuZscqZiSdVXPHJukCrNlroPo7dK
b7tV2Qe1mzDCTgewblVbqQsZK6+/Z7cC/2bXPrhnGmIjgb4ZT6VaforjrVdsE68p
fTjcgcogkPzfGrT2mz/iK6ndow1MVJB2JhqhvXbnVpqj2mABnVzkMKVs2XjPjKPW
0stSXiPU6Xq0XNAQRMcigs5AwtPghXq+hd6ws/zQK1+sLQOU587xDeIGK12W4RH1
IWO/iujCi1vu0ODRd51r1JxSR0PmjcY5XAQEyJlV7Zm5WvjOxmDLnHB/mWCW6t7+
dPc38RI7xHENycc8zoEDE3bKzfF/dHtssKJPwpXGwu+f93oPv9W0x84p1LVE/Y47
+ZIEHaxRaWawxJGc8T8FZbS0JPEoko5V0WRRZBDUptS+88C4Og6Z7mjtaY4YrI2h
DgRMi7fHX6iyqpCk50MkU7oF8LYy67VKa5VyTtMKYlm9c84TaQmUEWfg2lHhpg5J
331s/f68TDYNGn/bor8GNzLHJNlVp+oKz7U4lVB9Q9kGyOzy3InmJL362u/wtuhh
ljOkk4mf1ZmxG6YdfHnehexUP9AzZHjuBrI0jWemve22EfTfnO8PiOjdHOlvz/aa
+hyxrUyJ5tmZlYvhxSlmjjUZ0LJL89q/mMR4ezb9eBB6lzJDBmS3tyKUck2fvLz9
619803qDcOTS3LJtj311BgsvlQ2YfCHfWQTOf/bBRDpIM60YYGPkfjcqljtWgsT/
21kGyH2o5BYmpbvqeYr85iqpGeiYtHssrjyNs65/lBcDTmPHy7T4OQe5mmQvmVs+
fm/owXNvarmwVOBOMgvo4uC1GE4dK01ImwtxxLIHoTdx4szuw3FPB1gVr7CBMwtn
n/qtv2KuuSxs4QrGRxK8XwCpywLmIjEWjoAJ/+iKwNot1kqGnbMRMbMMQ1SWlPkx
N7PYTvvuTMrAXLZW3/H1erp3Iqp8+7L3VtTvo+j3mnhuL8TXNaWA/BG14WiOwu0T
cZYWRrPOtibqZ/nC/3P+vfGDGnxZT2zGVF1T21nle9geKxClIru5FgvwtOu8wNJO
0k6fJ3JLbQACGceJGeU1N9s3OwoRyXUs+ahjXpVbpBF/+ja5yiSZPUrU/gnHR9Wq
5RpDWaWX46Vg9Jo/UnQsILi2or40Sr6WFLSVl9l9Qm4RYjbZiJpXATBjEPPgrws3
JnHDtD0ok551ci2fl2yAP8+hu4DEL1GJSesSBdPY012mGknGMsy4KeObyLCp8oi5
Jk3peeJ3tMqJwLUE/tGwkD/LbYfFfiWJgb6QC+JdlC6fy0aMJkOIkFMKPwUp8YzG
tvDzBCNiQvntLnqEe8+MWkHSa8EL4dXpHb17McnR498/uXB/hbD/sqJW2tBt2yEj
AcIbGCbjAgNYwfL7bpVMu/KP8A0pBKoIneG/ZYIlr04DTCY4z9lET/W3u3ddlA2A
gLzxSoftsMDBD0NneAvEhNp3pwMzTzXqH7YuR4oOgBa+6CAK8p0fE/T3bM/7oAq9
qhCa+MH62Qz3h5BD5g7cgvtJLBQYFNDj85fnyyYW6zU1OEWiktIJ1HEEzVwWRK7A
Xkiny2jYVMiMapNIFMB7cE70Hhjol6F38EDE+b/MKNaZM9DF+Ql9dF42FYl7aWzj
7AH8FjV7ET/Sn+vAK61YOLuUUgQQFCPwSeXFSQf22GJcGkkMe4ni9ZZEu4+GILJ7
f1nnH8byAGlvhWR6yK0/KvIq+Y1hatHhK+fVmS7p0pq23mqT5xekgEVa0TN7jVW2
N67QkDv4K8OnXMjjgye5iOS5h7RzxzEPlMC22+sgN5Abaiw0ekV+FTBhXOSfC0kp
EZ77lKsu/q0dcmLjBLZTx54epQoq1T2gLA3jHFmgv5DKmakfwJF9dz7WcUTM7cqB
ie9qoyMtkN4WReALQQegqJVrD7EdjQoVBP6RZ/VgTzT5E9nQ40+jfmrp4kRGVr69
ipmWxgCbaYIcFe+8QS6dqYflkE2cDM8umluhOAbQzhslo2t2cO1eLE3wXtlnZ2/p
GZHwKQkDmPTYg81F6L+IU6Mo1+PHK9lQL8YTA0HhBJYvqVyYVQobnKL5zV3SmlIO
MNK9ZKm/L+ut5DCxosRynb8BG4bJ2qX4AA2yOQxgZBcY6WXfr1ZuQeE2CH8JlxzR
gYLwDUK/D9IOjXs4/NloedXDbZOiVIkr0lGrZFK0htLEJ3Cv2++o5R2lK9T5Qiym
MYetj+I6X8+VsHpRCLsubL6RCE1j29hEOktswI1/kXwOiH8t3ritJWZlwfpDXD8v
+32Nd8O7lOLsVETwqz+RSXYn7cEkrM8yZD/JnLzPyuSWZkjpIHQFQTN5EQJPM6oZ
URU4zqlriydJzsIFTA/4wydLCj5ho7CxcrrJh+pqkBSfvfLv+U1uNBJdoKaVCqBv
gSLUXNuFGK/DJ3m3Nd13vKPV4IjMvpVcUhukFIID0Zg+jjaXwZK3oTcceGtbxs7Q
1Dgtg/a3EzTMWJhpn8zW/fTOfKXHPxWhJWgATgP8+tc/nd+qThDyoM3K02uES+HL
zS81f/9qiY1sgYy6PjrS2dbL74c1D31qAiPTovszInF3vbrYX4u1fOL6epUgxzE0
aM7KhjmDd+RLVFypgUZ1b8h7ICxGfKc94etYl/EnDdvqNsKzHrvki32U75J9fZR4
oiNS9jZlij014mQOg9R85+ExQvbFQ1gNw2vyK7ZUcLyjS27TfGIASddg3KOL3VTD
xF/u93cxGw2BV9n/rNh1PQmwqVWhatGmmmgx6HYQBOok+IDuchbaf+Jrg/zzog/0
G3FRJ/bSLNUDxwNt2pMSHba2E1fqp9N7sEl4E1v0T3ERclYEK1PRAVqsEC38PfwX
HVLH/kb5mZhoVPtHAHpojAHTD3bijg0rnssFQy3gvgb5/FTvuyVqk0AzgOFnIAr3
DF8Hxhr3POZMMefavnw4z9RPN4sjsznVATQ1HMg9kLHQNWZSdAIfhHWVOsckaCAX
nTngkrYqYuIFZidXRW1gcnOAEWi0AgBhUj4K/j4pXN4sMwWun2gy4ITx+S8FGBX8
WvywpHn9BPqJCO5idK8YN6y1DgYkqB7j2uDVYBreyfrM/+ijDtnHK3EdsoP2psj0
Tuce9QFh29S90uMUUtXiFjLICNjZhhE1l4Nl2dJoy/YyJtjEkx0HOOlFe/DcgwBt
FXEw7L/J0e397xydhERDBUeSUOj8wkDKBEJQZWMoX2tuFkz03VonGVVuElY4OqoZ
+fYRxgi1J5SvqSUSd8Y1+ZUEBhe+a4oMLI6/FIqmh7cQRSl2q+a7HNPK7SuqVZGy
if6whZyOH7LD3tM8dzt+YYIV8LOdlo0VVw5E0jCnbaIOaAKTOx/ulTcNTRB0/6fj
pnC80P7bk9iSi7wPs7v/PSgV/h+TNZ1iDAHxh1FuCWybvyxBXXKwzUblgbjk+AVC
HR2K7aanABCJZGtjGaPRmYxIP4q6VkAPXUsyacYLwDUU86Udr4Bxmc7eG3sRWuzC
VF3s93xWL1ohS9azSX23aW6uDmQtcbnTxj9gdjWGPm30LnLQNQegJky9L1TwdPeB
tCpWSrMmzqRiymXcl13qhQvExfCJ7mXzwKbI3ebq+OhZentuJbxwbn92hZ3JErbh
B9Fl8pShT9buSgoYu63lTSOgJ54VEOQ2O185C5j9PGfRwY9+r5naXq6WRB89NHJO
KQCyEOnMi58XPhkfPackkqegW0UHP+BU/Vlr1tT6vKsnGoqHqtRdMQCCp62LK5py
VLvZijqp/HU4AwAtqreZono20HTt2t7OtXrVeiY0Guco4bs9BEl0C/qI3xMoQHv+
EBV9yX2hkXWups/CIvOrBDcZkh1ct486Yw9vx94bak2cirh86crD0tv1r0TpEuhu
0587eFPWyFgSir1+QmkyD6NkcGgP5IwTiCv4CJJZ+ZDqiHhauMC2pwkmIB9n7s2K
CkBKHFbn4qW5oRjnUfzAdotUrQfgbDZIPRgYjVZJo1D+h2aUBjx97vgxFF2VcU+i
TGIRtQ7lpqb8LGJsq0sWMUmTyhBX1KQdPgVbvPq7hj/iyiOz6sI+BX8JQrU6Oq3g
rAZstw9hwV1oTQpPL1AWNLLJ5dBEkmdJZ+bd1kfptCsjzOuqhBy4EZHvXoHXaOWp
GCNtpuJ5ENeU4Y6V+CVMuzSwuaglUYD9s39eGO5sDDVZ3crO6lkZ1sO01cfjtdwO
ngevgn1Q8bJoMPe02H2qNjSuNQEPdAFbhLNngOB6B4L3Wt8uvCHXtu3ECG1mWsGD
Bpd7yusxAVnDJTTe1opYmEP7QK0U7mCMpOiGsg3frIWG0YzKd8HkItJJtlERDG8V
Gw3upmu2/Dsi3z65Aq9bymsptNsfwAsFzpezfaniM9spReUXqSSCeEymmOUBcywy
m1nGdY55GCXFIWsOTWFJ4SU4axZT2WjWrp7xP5ZestpNEWH1YfEm8oLUUVeY4kKc
37IasNWWJ+AuH//uqp5bE31+AGpg2UA9wp1dh9JExOkxXSCdPXpiPdPjkIEFoZ2B
Y9vB6UFqGGuy8SeZAlVlfRWS98D6wDfMLxvgnjqhVTmgS1FPQTJSBR92VXjr+42L
2Qo7lDiX65pR+31kwUKhRexqxlRuewrlYR+XPirLAtknWfMGhlubpXWql7+ITAAb
hklQF5yCFv6TXEcrYjQZGNXKZOc92cn4eD6LLq5jXKvQzANfAfvL1wgSUAay+qS2
TQ5jr3hTJEGUmwSxGE+3BY7f8V3SbCHW6ztj5zWiddWn4v6uYf8uAqJYPxC6d7hM
3qMS7Cq990l+Y76oQoVj+6AS9Z223+JWv0ysYO8fRZkbjNnuiJsgu4wFxRz6tZw2
WQ6/Iv1lDk0p/vgldPmPS0qUPkCxdK44pVzIPABd+ZbM7VEsU/mWaIxrMkq6B/Ow
6dzIhWMe9d6lzOB0zNmg7uMrZ7uOYx4dQqrinb/xvWnUqL7API/ciOesYvZXgOAF
l2OZZ2ZsLkXki3j2/s2cJrD6CTI891XT30MsKd76qsiJaOeZOZiltH3JuknBwLHH
xUC1C5TiNchkSWBTmUOlqUeHLQG5KXRysSwnWcUtJr/UrH4aoKzbC81iQ1d2NCNX
Ak11fHKsCr7e8IIJUr+p/6sWyvIiEXHOuktAiWHD3CHr4795ydQOCvT3jnoV9y9Y
nx8Bt1E0iOAPUWH1nz3ijUKv6SpvpgiZ8PUWKQlX+bQs0YlKGdEyZqM2frnG166J
6UrVaeZNEFp61GuQTjPuNP0zmGeXpU/MuCh2WHgHb2cnDRelLSkvqrZdFXcbRren
LxZAHA5iLrifFDMgOp+bzzgy1d04gGWp/ZNJ759uL1imSulhbscMxJ892imYGsyM
w1mncYI9ZyR+mG1WSe4EXf8SIiaxFSgW+/HUQQZn4YOzDf9SbuBZVRIZEAQCmVLp
W+KmxnYDAdOZJ6SuKGhnzkLmuZJFTY36b2EMszwRLemwB90TL77E9Imc0mZ2EIPb
rKp0VeJcd8WJLpP/LHRl1qXHtlQFjIBLrPAO0Y7kUfr4mTYJU16TmTyblfmqXbtq
8GQIILYdMRf2JdLDRWaBdzx8X9HCdXjGsV8Y+lySvdoLsm3o+LotT+xdQoJ2/M/H
XcArbIeFT1zdNlGFnQDf5pvvY8N0QIITGpYuRU88lZo6u3LTPV7Y/34YlL3GUVZB
aMrjxsP+8MNKV+Ltp8vYtlnew8ER6Wmiq4nc1EcN2tuGWAKfVbDcbY3Ts5mQ4818
VlV0QF94fBHMOOVtv7tJSgfpjBpoHgp9yTFRHkJ2YyynvcqeF7f+2TcGmrCkZNaj
Y45VkGQLckXPwvTj0mDJ+NW6rt3WxhOsJVAtQXgahze8uM4LQhKwVnJJxHuE3n3Y
53ATbJ5kPi8gLFAOPQaLJGnZ6leyjEe2yvhRJn502rg7DIGckv8cbrkUAFov9iWU
k+sG6bDHoyFwQ1sDRbx0Aup3s8OB+I2xSl62HwCVKOq3INAux4AQQ/gG6C5VnuJN
p6x4DOKhoKxaonj3QwukM7ryIiB3WNGxIJOTvDTPbSgX8AXLh4QlDMR5WO2Aw5Ff
7rQcR7W5K1DiV/BlJNQRZIsTQ9vHzLpibtt0jO64vu3lyOBDroAh0k8KVfQ+cbGc
IfsaRhIqaJfd/WEqpPKuzcXhc6G/zGjtqIndrCpcxFxA91HSyZWovmrx1PW3jSkn
jw+FXeSSk53gxxu4PfklHKlKJKQgHWBzu4DavfWM7cO/EGwrnUIyi+QhFqoY70L4
PPAb24dmznP8g9FrUGvASDtyvJWifyDp0D5F66WTSDwGrzwXzfstZVhnjXwv+d5C
W+FMeFD1JlIkVW67St8+8RrZoeU5wBT48SDpqUv7ceAW8ITyzHubVb0G50A7V9sf
6cQsP84lAlEFfQ+V2rFSlRzOyIBYiO4hmvopC0FGtdwbu0Dds1/ZiR9w6aWqAqFB
maeqmA8FSvSW/ptn9OqSN3yEyjHdl46leLbUr3RyQePKx6uJ59+YvibtgBsKXYFO
nirAhkzwnmD9cPRBgJn4YC+PvAidKC4bUoBLTJ4ot+YotJ8CGqN46BfE5DpiXezx
GvxnqdPgk4kUYhjC9eCo5OLG3q8HZsF9KM0H0z3D4TuJoPB7UWfUn8CX111PEJB3
utJk7gVMkR11X+S99Q/JD/Y1uQnTLSEf6boU5mC4ain6uycfmCABAotT6EV6Tpq4
tA8Uf9SWuuP+ehHgZLkXgdsPI/xlRlbv0QLRffyMDWrHmMpM9WN2ot5TNQtc9hFt
/iVab8PzMZYgu1izp28fb62Yz0xER2Ks1/sFIGZHi9brJEVO2lJFZpX/4z7+3aIG
cqctlr22slcV+/W5JbfhVat9pb+LTL7WtLrQJes9tnTWrHT9kMUv03KT6gKDqB7E
Jeh3deZyM/3gX5WZ9dX98dehlDHGB3e3ZdecgOWQeEbVQw+4RWvKNEk2lptjDXXM
Lj6iZ6IhXUCYkYX8v+Uar/a3xaUjrUSM26l3Eat6Chqwircx2EvAFUFNYTuxjWL8
MIywFiozsfwtU3bCJ/lV8Do7IJLJSxSA5M7kDdrOijNLTP+piy5atKKdM1EuWCuw
9D5QhRhkGFYzveeDugVoLVgbdLNtOSE/ALqvLRvcDJtQ8+Usge7F4X7K2konBXaQ
e4a3Ea4mTwHyzYTFOJV6CxbjqvYCF9CFP1I0lIRFeNNNpymVLULgve0PTL78ApbA
12N34P2rYjjUFNG+hBJccqlpnMAgwRpFEyT03kDzmDZLBpTFCyfaplSPRwvn75th
nfREQcrpuTvozKVLLwDbn29qUnpJWAIS7ADj2+3t3go1+6TvZXG1cCsjtEovT+Z5
3lAH3Ked3PWkFdS2f4GEfylPISlU/9t6mmAE+DJGK4Eexb2/J2z/eFp095f9U1uT
ZlYu+7+fXrV0thZ0B65HgDg68B3ynJGbiaLUl5ZkxVSxrp9Ff5Lu28ARso8niYMC
pC/+akEj1fnLN9LzE6p2MhrcG0mEmFpnsjzDFHgrUWhz8mu3MkBTiMfwW+rhVcVF
W9TYgupqc0Lre+YlYjoB5EYOFiv7rdq+nuy/H4kmNOkUOH8IMiP9/q/usfpMLG3Q
KgfM4ukXNcJdQqQefvBJ4YgD9qNcQaA8TPtgCGCKzTJc7TZZGgNKR5DWi166NepC
vINsNETLt8x0uLGPFsegVYtvYkk86wiy+JwH02E8A0boT7RJDpSdmu16Hs1HRrQk
ZqNVuQ8szvTXb9hsJ09iAosP6lMTw+pdL7TxSWX2xBCE5jtxSPvnyYWEsLWyLz5+
t/ZTIc3Z6X4mNidKerD0IWv2sTVjCkSat7ygx2407SOrFABenJaW+xuHOMq7TCUD
Lg/TzICoDaYQRS7Gh5PZzxIaiPetnPFowCfQiRaSJ5gwJj8bkUKZdLRv77tkRcy0
xJfHeCwBic7ALUpsi90aYOOSYM1V7mCtssTiVGb+v7/f0vBwgCsM1E+59RgY8UpT
My66BrBqN7yvrqgJ9SU7HREsqKJ8DRzNtGg2xVIOh2A7bstu1OP4pP/n3p0SCylo
V2tJqwfHvYdvh91lS3EDWffelIb6nLqZwGJT10sz6kI63f/+XShp2KAS2q6SJOcD
cyL3k4ky+4+jer6KWk59aZruvRATdjsRTO/iMaVWwyB2+2/2sswgZjT7kvd9COv6
OR+jqAini3GHZuufU7Iyd7Sm1unslwYo+Awhg1X7UXn4owl/mYwkiDXmb9hGnu/p
GnmOhavjQw1Bslf5geb8zs7o2Nq+jNjvRg0EZV51AdhsM3V8lJzQEyf4bzrjI+CU
7RUZMOKE7zPUqeGRrG5/Ah9fkFWXbQtZlzwG+pRfrvGXH9nacCvZdb22mYLMoJTL
6OAplstQB4sIHszgIzlrTLAGlHAKBzIpZH2oz4KhVPNLrJuxZA3CKMMAj2p/wf9x
OLZ9CBBRYVkgvDRkYDIJ2W/kFHinxh/iE1jcHosNSD3RlqYGoUtZxw73HIkuDbzM
tKrlkUv7spuDpzdJ1yisjQtAQ2WZ3kfNhcnyB/Z5hsTEoMiuKmyKamu+Pi/AxkUF
gPtXm8BgrI9fKTgqflXgUZ+ITGJYbJ7HL7YWARD5v2JMf3YxoVx9HSwWFcz12GX8
BzPQEbwhXp1l69S6pglKm//whXxka9JfHTGxDzVZodrgQPia+xghR2VJtpft/56W
13/YDf5WS9Yz5h9FuOTp9FO3AjbESvUNwwdbiFj2CmVhhDPaVaOPvm7GgX+5jAz6
IheOo6ggQuFqq4G9rRUwbMrVG3RRkGK80CORoHP8ODfS/2YtyxKoB2pADk5hcmsb
XCNy7EgegsGQ8Mk8zLpbi3xvUOa2ixCpMKyznrsDU0A2KknvaTh3KbM/CJyOByh9
8Dky62J5FjDIad4iD26GKaD8ZDVn5mJjSTp+90enbmA5zVfhNpprNNWRYq1DnpaC
am1Gc8wpqElIMatj5CFXWxoT6d98uayuhQw66EZYQc9Bl6S0LiKP1byGXb1gJ+dh
qPiTo9Qb1ntqIx2TGQmhI8TxYpq9TCgAEz5vl6BdXhqHFH2KMevhI6u0YFY/p1FA
YS/ctfAwuQRS5J2sVtLzLpFB3bq0ofNZY3X6lwWP4IPpPg0GOpm75GeT2vDpB/Os
xkH6ydypOweIh8EG2UzPy1VF7J8eaU+fdcUm1lso+ZAk7150WTFIFAUJg/heuW36
ba4JhbCCIEv6bymIzKFmbM1c9Yj/qa6zM8HhrDwAvuM62El+VN3HJuD/4+i5uKV+
F77EZzxuXeZOEiErljQv+c+dwXrYAXQbdsbSuqxW8O5/XNstsWvL4KnYt7z6jGFM
P4KmqIOLe3sDmgLZCOwvCFPVFUzRn7RU7fXfjG77p4lWnEyiUCipu4M5G9Nosgqb
By7D/abADhNdb2oyxlHJbl7U34JsUAdFItv8z2EvqZjNCkTvv5x8kHMwoZQOYVfW
zfXxPRiaNHT+sHsm3ENuiMvtkd9efTdCuVc6l7qR/JfnnWxwqRSdbgb7U4hU6xKy
FtYh4/+/21CBbP4RJhOWwk2WkeBQMokUV8HNyRMlC9dNTt3MvBcFt0LOpeEjMOCH
djgdOayi+iO0RxsaS2tLoyy6FgjWT/VwTw9aF8tdSoe0BD8uOXupEQiegueOBl2T
qERrR5g9DZgH8+GVm0pAOBuK66/qe/OCjTmtNFwK4MFYTCp5SOA0wBHBfXUc17J5
0InLVp1zLv7oEeeII8HTFRX1DcyqTV2QjWgokBahvHxrGZv923UQZQJIH9Gdvj21
x4BcNyuoXI+7CrtaAfFPL5HsQpfZDUEbnBm17YofCWClRgkHaYK8JeDp+Vp/1vu/
vd1jHOs9+QqbTDGBDWQv26F00oNRlW3nuhAXVD2p2b6gaf3lP3yaJU8dkfGF+YaV
BspUcdebl3KwhfllNZU7CD5aDDIxGULUzaVrN81YkT+opIanuuzy7xc43dxMr9NF
YScOG0TmqBq97krGg3a/YI6vGbRc+1RBdawwx4a+XChaNmnJlTL0Zy2xF6v+b4oB
TweZ9Emy+AX1/jz6X4H1h6JcyqFiO9bUeu9P1Aa6QeVOxS//HpOTVOyQU+Z4Blqn
/SHaibW69ZF6z0dLPVW5tW7Pt/X2yxIJcbEy4OiFoYOThdfuJ+4D2cwEfTcBt4My
VT6EE0q0MgPPbYGbHQ/W2H+LDcoCMWVrZUP64LlM6sJnym+sohcf9kwFEeHKXLn/
amc/b3lZRZDVcfhI4ACd44SZIw6EcEF3sYu87aY1RUlp1lNkX9lnsVeXyqrt6LYz
DbJC/+kzCVnVmF/soYaD4TYArzsL9OktyUgEJiWhrYrqdmpGpw9pJ9h/Q43gHJmi
CVkPWmHrlrEg91qrVSQW8h+5VgB0R+uNc032u9EAPpv3y6trmW1XSI9HgIHPv13K
JWVD25wLSmy5pAuEUSOJ73P5YpuJp3V/kDcXsMtv1fPJdMxbnLBd6nADJ4wFKAZz
J3LR/0Ora3ZhvjsK4Z/R096BpUcyKBDxHIoIiUYX4r3mRVgz+aDK7j55FsV0dm8Z
Ka/WJpJ8iosNqZMI2Lrz/Bj59JVzMdCRE7BCBjRPSkQqm22k9+nyGg18s1sc/wXf
ZKGe7ssv7JSqf7GM2dXJHsbQLYx/A/va0gd1iHqpoK6oX8/lf11tiIiSzIlHT01/
qsVK/zPpBb/xtTbANb5jQXu/0PuxZ+I92knZQ4Ef3Gwnt/4sZlaOt9dqVXXptF5/
Z1Dh78cDC5R5+MH+W3BmmFWqzMI8hwBwDzBwq7oMGUjzeH4y0GbcSjwZPiVXUAxS
KHqd5Kg5qIlmwFo0Q3NkgmLOt5Lzs9tio1OD7tZwG3xeEKc3TM9PuUNT+CQG3gcA
iWqboD45i+/3Gx4L4OggURtu68mWrFL2vGqyhUl6zAo+WIYomIruxs6Htklv3qen
YksGOqhSoZggMWvuW4GKpbg7vaxyQGO6CR1Vb/9D0HVHp7MdTZGDGUBTsuq8ygG7
ysj60bzaY7M7w76jWNecOYmut59k/LLTEHaU+XH4KxmwlU1CdJPZxZzkiRWWC7oe
2zJ30Zf9zFg5WixTtEQUu9YgPG6/6+2eadOQCbrlwC1QA2XowJYmp4pfutI6p3TO
pF5k66K/vEjhdhO5N9ASZl3+VAoCxMSLR2VSYLPZqUxu4Z/J7iBREQdV4T7NE8v/
6yTIZ99xIixcqSMGKfZYMK929dDpp8b+L3gp6tg1rex4StFH5hePEM1iMpseHxDJ
oDemzu/+UJOKVwzC0ORgTHE2wASANPoR2XPbEL/sIBgSna6LcpLC7Ck14ojb72ag
XNrC8o61ps9RWdSHFHrS9spvRcWn09baOY1CphQBsCKwQp+KgeH/ftHDN+CsSqAI
tIkndp+zj1CJ9coUR9ukVnW8V8Mf54JYDnc1aII0k2WdzDb3IcuRSAuXpP9bCMVH
pke8OzRW1VGJXA9waf5/2zoHwtHlQR1EmvdbyA2/LfAby1VAbAAP3ItWVBFVc4wH
Hlh3OCZ+nF5EmffMzh6NJBCt1jh3+g6WdjMzZCjOXQFY3pFCPz/eTVYzOFPa+yUH
1b13Wp4IF7cSphGE1MuayEmfdXq+HqtMt+/4/VCbQM4+T7okeZ8AikReZT2jmdgz
7vJOmOHuxb5tYrbbHrA528Nv1EPtX/gOdGH2x0e14yBaawu6PU07oz7NvVOqBtsx
SXgsP39S+WSIFkUe7sNSSb3k5U0H1ul+K9HeQeMhzCBccpDnm1GYr+Yd1yO3069v
jKvOOiteqNsGto444kRqqdjKZnpOFpwz/gtL04ZrFbRKW8tOj0tnUAFUlU95q2Bp
z1UawWRdMNV47hDQ1HCoO9seXTGWp/1KN2N4JrVqJMKN8AUyRfAUhjAkUCtqC73J
Mf9gfVxCW53nvFUWO9C3qjRm2m7doURXoMjUOSMSr71P8gAa4GNI6pqt/X1L+ygD
fnpSAwJGhmn7Uujuja6qs1bKCUsofOUhFbT0M2NaNoQ4xAUW8vF7Tn04UoNSpfx8
abZ/HW5evp8sxBMGrw00AzEHezbXr5POB3VHwLkDpk7Tr9yZeputHTwMi0s22S8r
wCLthpvfNV9oRX0LQbmPa6Bd7loo0YWR9F6RjHi/f3NjxjJa3NfnIHebnfo8rX4g
2pFAX68NnqBX0lB3Td6tJa30OvOW2OfkHKSMECgVa9UBGqbqaeOzbyG+48bAsPMh
6JpGKTjaq1b0PuvkTBjk+czn5cm2bRYwGMGvOzMuVi+WVlg/v2tjDd/kp5i8R+nG
4uwLp4Lc8BNLTzgR+1ydRKH6D2/SKXBEVDpGKD6TmvrUNfE2P7FUz7i6oGS88xjz
sqUFVveSDNDkgqyh2WIgeyq+adnSxSnpRcCKJT52biPdfHrqCqGfgxT60C5/bvL8
aTQ+YxWNstVwSQwVB+vmWeCXu65udxlr4a+ZSvqgq9wi8ZSVS3g3l5qjlZT0D4cg
nkTfRFbf+6uq7L/V9FKnNnT82CbXS/X3fBKdtH9C2jkCuT8+xpBcvvvNdIJHnV3k
FZ9VnTvoGbzqddLlR/pB6hILjoLCC/JvhbAatdW8nx2QLVLPBiUcaav+/gycHvoz
7QOAWS39Zegl9eCo9rIJuTjb9p2538AmnuNfWwGGTEagWJIgWfChW5kE+Lmxw8Vg
g+4X11EIk+W+A/d2X5o01YjOFY4fz+miu0gce7CS+Rr1XkqM7hmU1OEMDdflSJlO
QgddvGwKuXxIP52fbyNrMco0kHw5IbbQ1twv4lQSHfm219Y9Pd6nY+ZYmnXXyIln
lnHslZQy8CUYHkpdo0cTf6zps/43OGegNmiSfL57qvSHpvsyHVGnhEBVLkAOGMOl
QKppCqT92OaZl5VeOmcbwiD1Gsk0oKv9bVy139B4gBnMt7VSSRAdpborOnC37D71
K2Dvw1gz4AqmdG9UD1wJzgC3MR+ORlDpchqjtQzwKoYEKSHXn360SUrzdcNMtmYD
rwEBnJMd4fkRO9LlUCtkPaKqAMkrgKmVm0W0wD6T+KZpa0UY0tGuaoY23ymOX0su
xt9c/YkJpTYcDGSJTgafmkbaiNXwC/1XyjmWxHmVF0gXEcpUZm/4pEB8Ezd9oXFS
IgSzmZnLMDFP8Nuw2CYn4DiGe0d+ChqMibNwjVkWPKdfvzjSGbKBCdJ1DyzkUclj
+Lsmx2rl9c8FLG9TzLV5eI2vFrxT0N9777nhUHjrzvvjKHyFhU9u6d8wA3Cosuiq
KmytkO9vNaxz0g/ynTdS/c1KoY0kfjDMt0+cHnCp+ZXDpTRM/XV3cYr2eVAchT+c
GmbZcCiyafZifLLQkCNKHgJgUssnOvH7ft07XpUZA7bjPDopcEXkF1ljn/ARdf2F
PbA9APj/y2zlM8xq4SwzcTh3EmgRq87na9HtUfo75vVZ0uJA7lQ54bXO7OvO8fqS
RADLfalkaSCOHTnozokO9JYh/u34uAp2BKmimxaRGerHIq34Gf3rCdPMoGNxaCHy
U4mFrGYyHrin8V/nHvBGHEEPY9WXZu1PJtDxKR6ecPiUrtCpc/DdUcQZf/Kyceqg
viHkp3fjAAsegY1L1elT9+P/HaMsGRzbmVEW/8b5Qr9L8cEDBzX3MqbXriq/evNi
d5xnVoF0fpGecelfxIomCebgH230r0MrI8Vn5+r+VrJAdI/CqMYMufr5utNIHdpG
XNq3yQH8IDc+sx1dd50vlCEbWBweDrR1nkx9vvVYkno38kdkH1EjdFvjS9JVlnoc
/ZvR+bgZNNcvYRym8PpDqpJOpdqspDdmcOo52xTA106otxRgtopBwxulilmkawvV
q39+wCC0QlIZ9ce5ukf2teu7T5+D5uotl3MkoX+g1mK9JY6HX44IPAiJFS0qsJp3
9JSLAehutyytxH03Sw3+oD/7LXBrCV3Yo6PeZRT36y/iVpc8XLJvNqMVPDuvZBw3
smleTu1R9FvS9VuT3YxRb420SHqq+/xFNZAEUz/guuzY1siKzlqpc9QOynj2ODyz
nmLhCp0kIwAl9V1PSVznAU32SKuMZReJQt+LPTbnfDIkqBO9YFTuWHIH/BoYMhWC
YvZqWcxT+11fg8On2WBfSR0JKopjxQwcFViHDgfaRHTNIJkVEFG9Z9P0NTKz6wVY
AqVgWhLgKiWBa8UjERT/LDJr6L9HwupY4w7leeVEbi1/28lMu2asSo4zbERlBk1A
1iAmJtJZ9KKKP8pVlpvjdvfbjC2vbc3u9Eae3dqzHATbcRkHBPaKlWygWyZL0teq
a3Yy9pLYEaiLbcQZRZEYqpZ4NlVT1KbLT1FJDEpzZuGctqIFYT1f718LgYkop7t1
Kmvfwbuxc+SH1Ts3M+MXAWbS0oKiATZA0W8TBjDE1R/qog1Ia9GBp2lpvOKtpVIj
hzit3COvygwAXhpoKlarFcOyeCNjQOTbG69hMqMGQe0ndHs/dAMMIHtW9FE2ShDA
u9CieZWukiqxRsK9e42WlFh3w9PgHvSMVxriqTShb6LfU45HiZQGPSeY0OT3bf9a
zr25nanUx6b3bXAUkJH+ClC9QJ/5F6MjG+r6UVvAl3AAitGVrIJs5cL5MPt9cA/4
gMLxI87X9j5934AE8PnKQZYbW68jRV5r+mqqgaly9886VSar5/38dEsd8YJvJDI8
8PXlEhBMNxG1vxPAeqm1gz6GrNrxwwvauENOOQdfDD2+9M87FyerhiMZGwt7AewV
ohYdsUXxpkmJlFzrQZyBcoC4/xwyQql+o5ryo+78C8JXYxwftRoqjMDl0dgynyHS
FkY9kqd4PQXIphYVfHuVXHwrtLzd1KMEQF4ADzvKspbZ4G1gDGVE6VEBvWA7slYo
YRun+DeZDsSCqHvcy5fHjIYvWf97GnAyUN2duT3qYIVpx9J3X0bRMtGtIFqfnDXr
ua11NBDacdukc6E3h+S4VrH2zi6ctTu2t2k6WN6PdGzjR1D9f59ltozDQX19lrq/
n2mI8mdR4qtS9gcKqzqsbX/QLo9RMDE2n05XR6oq7F28uPbnHSvCE8hUJ41atAVP
XFcIKPS2Ok5YJwlr3AISHuImCOCAaV5xTo/2JrxX952QPtcr0A42yJPIQNnCMnFT
T8sID3vcHDGPEtmyC6vImmQxsPPfF+H2HIv8SmceNUQI1hz09ua9HqOP9gJxN8qj
tWIBkvBTuSOsyT9HjSs8cDf3yK5sMe+hSs8FpcmFYMB1GPRrpuiIb/1k1ozFbLF8
Nn6kS69mFArvHlS5bGMYshLH7wFZgiHszGu4beDLUKrS4Tmpzi5XTQYqCucwyLIt
uQ/K8b7rOTKwi/y/GEvNJDw3xBNmnxyHdD99EwPY1C7L58U7tSw4oFJrabjycBqr
DGIrS4rWF5jlTIRsVSoPqWQQLnsBBCDyBw0pU2nCGzacGIOxW8PdD19KNtxay4UZ
868p24lEZdzFZpktcPt87Oo6hQ/sb7SJvi3bJDgG+37fGnGCU0rFnK8fb+2XqjWT
ALVpwJwhrIsNrgkgXI6aZJlQ5YmtkHEiEzEhrns+GvO0OeDDbJmtU6HAsRlpIfXW
2RczDjguP1DKRiQbLJ+tJPaR/srogAZKymPbdQotKhq1SVMHeD9S4PZY5hSw/5ME
Bt2Qj9z9P8KWcGjufbecL8v5ILQxEZUzIE0EZc02jWngLnC6itDT3MJR1JoBxswH
KIZa2wnlLgX/fyZZ94oFQzzKGxBmqRffaOiqosp0J9yHH8W89PnN/vEwDPiAKTlK
YPVQbyWuTpRcH97ddVJuu0lO4lF16viUgyzzGZjiKs8jW4q/HdjJ1NxPiI7fASVK
qPquJFJ4HEbovdTYhDMZoDPm72iCClredAgofbhQ1oDBEoXzg7WGZykCyLgBiUpO
4RQtYHakB/nwSbU5oGiTM8zVvGOE4dxJVPofUzCJRvZHAxLUSJGdj+we2s/Fndjz
CX/DNdHGcm/dp99Sx2gZ66QWcEVSUuf0OzYP9dWAyxSs8tWr/4u24nAddRuRIwSD
2v0nrRvOlDO9KYNmRxyyeSf8PPdqfz3Iv9V25Yp2I5nHB0OjcW3JVz1uYEenGV2N
dnmp1tnfbxnGJbVrcEWjy/0sdYpSOFKcx3yqqJysBJy2DuTq6B3AXvvs6WmDeydm
SwD++2mzZqfcWRWoMQ9RJ3ksPx0QcIGpMZhiZBcDTKgvqQqnRvhGFKufxAI98GS2
sfTG1hWOFA+406JOr8GGcIWFD97DofKwjOasV/A7VHihOGJfaLzmpMvsshR0AKX4
6ZC5ZAjFeBYeoHkhjK/XkUvBifDTrby/8/pB1ZQ4iHDQ99dabyTioocCPkYpk7fV
0D9G/EhKeS9fWO+Qn5DrmrzJoK7klcu5W6jl7SJwdkvhElOMnNRAN7J74c4x4Xxg
Emmmz4jMFRyGsCmqOaYQpe2o68HKhycHSxGY9XaqW2HoU81bOKfhWZU2VH9LCj9S
8uqtSlfclIObCx6Ozule19LS1D5Z5aXoTOt5vhsaVGLhhTKCojDmy5BClcL2NL55
tO6dTvUEjBfXEF5mx7UdqRBY7etgBzGtXf8w7rrrGPVwawyU7VUeg3QZ8MtiO0ZJ
zOYJShuxNFctEcSOD3LEflIEgwAWS4jmxXO2JjzJo+flvXos+LbtjGIUiFtK1ySZ
nvFpBMXIpkin66JO+9RJfaOjAn0RWpZlbAANZu9mNRDSekoLO9/SXIEz96j9Gd4d
tqvrZii+UXISTAQAnJ680sH3zjgk847+plIxbbfiv+oPV7INSFDmjG5lq7LhJStu
sC4/heVEBoYJ//IT0FlzRYCjyux4/+pQVY8vyvr8W5o5mCy0QuWzD+qCMKPrRgVn
3IRJ5AG2FkCLQT5RHQMGQEOklhjT5H43wDSEtpLhymNuzb9lMaQ58WcCMxcftrlN
+bxAEsBp5fG5ZkLR37EhHH2X/p4y9r8i9L7zySf1xOU39iFWqPN/K5hgW2EWn2+D
pvU4Du7GtcthjKhs1NZz3E/6glipxQW3MZSJfes6Jq5oZrj6HzmVWDyQaXNeugsW
sJP0/HKJRD4G34OmBGcizQvURKq2jPUAfuvX0TQgv6B7nE2uFEBJk424B7/suRBJ
TfpNIWDWA755G6lVpXY3ovoZ4SaIw3a0gl4dWgbPVzMtVbyCjK587SGCKhAip8sm
H6hTcPa+eObbsH/745ZlYRi2M1KrgsTKaDpik3xHDP3UYjeplhgRokscFhLSS6EB
iK/PsqV3IDRLs3s2g8Wop9TdvBeiVPR8Zt4sQE1HX/q4G+WWee22VdUeBvY0banw
wibT9yPxRB8pId2ykQwfQPWmoUTdl7KcIrbUZy76Z1K6lW7QFwCTlIBqkdgxAgLs
WLs8Ex4ElMQd05a9WwA/xDMBbm9yBL4VpGzDxKRXerkcNitV8yaqLnXeQhvIYriB
HuPlWipLQkys36CspASISOPtgiHd2ngiYQKLv1Nxdi3IoOsafE3VJdt8iPzrNAaf
uvFKM2c78jdZ1lRVhXt+5pUuYzwC6UJBrFReuHGq+7LwwRFGa7zQq9HLqyjUYrYV
zXrY4KY0G3TxgMTCTvg2ZLViDfwfQA0VLd3aqbj9IrMer0daaLS/+rCzhWnojCgB
wlgKnqqORVlMdEQ0QR09OncY/3CwvjvZTeiIg93P2ZrCG6HTrsQy5aS/sAGzZ15a
LZBJ0zySCStFweOWdqmzk0LWrSSD6h+dgVK/IR6uWtuEbbI6GFV9c1P50dzDo+sP
mo56awCfVdvE2EPa/wrFuR9TPl3OcElFbSowIgdej8AMEVDcAkC1FK1lJyGmw4JN
Nh5gHzUIdtWfT4R3KIxDOPn2chTxu6EjgsHrtkY61paVXvSXenthQXy52jyWiXNX
X7UYYHXG4QyPb7Tk36d7sX7hkzXxxzU7AAg1Qdl4lsKPHS7QAmEvv1I64z6Piwir
E1AWok2+pU429jAAtAUNV9hEQYLk6Z5pd9xMHwE3d7Gxmea1/lyOHKyfPvJtMTyl
6FoncKD3oO7Gvn7pyrv6Mn+5UN6oj0AZpjKTxhVGZAggN7rO8YUzHIuxlvFwdcqg
8PNyfqW3STkydp2aFiyp99XGEBKCYN1LRx2N+SHYrXPpNaGLJoKu8AVizOtOXoSO
om+qhzZEKbYzCJ+tCOXlS/jT8rp8jcTzel86iEvv+1S/nA/6raMghrPu1Dxikuug
YRCpToKXwxoVshnlqNqh8rOeYNTRtjxo7Nqfm3Vcb0BcZWDsmuiU0x0+8vbIQr7H
Jf6N2vvPS8lVYJgryKJSUf/jwKpDgEGlAVBe2+A1dELYrzEF2ea0gBryaChc7xU6
62zeWLdgI9QKpjvfbJCZ1aEo85LWdI8e/dY0S9fGckM16eJtuxDIV3K0tguTHhq0
0+9blJSl8q4ot+UQQwWwUoSW4rKgP0jeUupFsOM0tTC8oKIobTPyQFpgkGYAMBC9
ahQHb6w7zlQOWnTYdcS9nNbGnS6xp1AYsD3q0uTSVjWA02qA6o4+uLdulGpOjzud
EXMq/91k4G7rZ7ezHiSACrLMIL4VN/3o1A6GS+FPalAFwrO3QeojWeIWuTkboQHp
7JFHg43i8mhQLRqc2k6IPhYovG8MTXBINCvDElnVo/AXnCnc0z/OQpTLI6AgiRKY
Z3+yLCqLxYI6UhlEHFfFuQIPADfGYnSIO7kB+vGxIWShdDeKvt/kuAo0/SqUaBIa
oLWga/NJ2RqZ3sG6pLw4tXO7QviqVDGzQmZU+EynJ9OGe9dwb/zM6/AlLB+ivtDV
MQ4BUDiy+IM40lWhRRYsDinD+6mllrrGICeea09r7gc7Wno2I0lANHmhixGMbs44
GuOiSuzAVJsrmgUH/b9GFd4aSt0w04Q5TPEz3SWBt83qyWxLEW+IC6IFuPDB1Kjs
Vf7aRpXwh1T8iJIpbeisJigW1HxJovj6J38u2ds5k4VaZ+2oZ3MtDzbTX4xhNwDa
5xFk8/i2ktOI7sRZwR3ncuprGuiadhYK8u8/1piEkooeV+xSfkjkWZVp1a+TnY8n
9/MlCddR9hMbf0vvaHZN4FHQPQ18ooe15WvwKf0GWHIHSkbQdzp8NyH5jrV6mxUL
TpX+NXPhBELQKEpdoPraWKH7UKvl860Pb2o6mJdfNmAadMGXXCie6c+CAiIqk/D5
hW+rAzXGrZjnQjG0mux4DbezqTkYAzQnyPpt8zO9DuOc6MSX+UZ8eecx6wYely52
ZscqreLSkM7GdqhzcrCznDzr55e3Bg1kVoo1JfGZOWocosfLx6YYripo36sC3Bpa
8DkdloOe4VpOrNsmz9Cf4MTnqmKtccW/2994B8xT+ta5seC/HS86u6Wf1AMl94ha
lCOUxkXWot0fT61IreqPBVtv9EM7qXasWLAh80abJALDt+IxBEqEp7oOVhXwAxuX
q53+her0nxODazCXYf+xIIRvijcGinkNHi1J3UCOcw4S/7EZVYR4ssToLwPPxn++
O4oAfKjPKIcdnan1z9OnjqgU+WtgPcEUDPpy/woNBPwkt8JtgxekER1uq8D6wNRe
mbW9+E+jN+nTman9yE/47aMukLAemmV6qYer2mlGj1dtZLkCb01i0hvz8/SNrV35
B5ot46ET1lMj53MN57hSJqw02LEfZYPEpICk3ryVtAPN5yOeVB39rSa5PFkzpLov
I+9Mx2ui77woPbHg3YWZpzN8569P2FLTlRHwxrDtNOKGwNv3sdGbMTFhS/F3gJxH
j2C2zore2UqImPhgkZoKxh5iPxpt7MxdBVCFGj14c0yNzT3Ka1R7lygtqu6yFF7T
cwk5FQWWbSlglsrJH5lXLqVEr9PlalZ5+Nli34RkGdn1ieVejuaq/3OxQuGjdGbf
+tfCdrXzffIuUyW7oR10VmH60gv4XdHMQGKYLnXsgPfPhOLsbD6jRrtorxfrdo46
RXetvmnU/MdVhWUVwkw7GmTbaqDnJyXa+4+QIgfgkX9js8dAqoaXwVKsnH9Lk5JT
W5NSCROx0nqoWvgA3GDbiF2Ud5ocNO1svL8oKI+aFEckS5dIWIQrLaQU+B/8Sftx
QT9kdho8h3AHFWRXLlfJZQUOFzYEp+xvchCtUq5h5qYiwK+w1oB2jN8j+t0Vsbdj
uTthCbYT2TzvLir9GnVRnnFHZ+ZYOoM303z/5DYPwJnZ9atez7Fc/t0pAoowL9ae
6WzBNnQoSKfE7/L4gx2ueH0tqNgPXZTHl+ekZXQpsQAjtpgz2lbaaZF4Cn5SBkpv
vE2+yUz7Cjlgq8V1aFrFvybyK3JVTxc35YiWxkhzyWi7kuCQ4IGSklJST6AphbTl
U+idshbhb1Sb21OuTSiDgHHxpjL1qOEMNIz9OKjKZIhZ1+cPIKv9b4vR8c8jLpCV
MiUH4iIEh5anFCWnOE+ibY8zelZ0ecm/7S5R0tA0JImUkPQUPtEDE3Uw9wlkZ8TC
miZlyaYZCuPjzK58jDKm5XP4kqqauXBGQsIeD+TSAerhykkfKSTae72A1RWpxD3G
dWaUC4NHjyC4ROqTzcMwPZ54H3hqfMYlxsf1O+D/VoggNIz+9wBs5MIR4DuGjUmo
ZRoAMVfJMbA9cJuj6VmaVabDeAIX5MR6slX11JHeMGn0QYZ7TcpRXrALorYhX5kF
pOC73F3vBM5Fzms8CL91KnZmggAroXq8A7HJbx8QAuq5jJYyalQ4PE51iVaslGfd
e5mHm1VKR6knylB71ZEbITHqTXqTFaWPfYEC2sXhKGCD9a7plAzvLU2cNawXUTJG
BlwHNAdR3ZTsZcNQjCunOvRwKAiDwG1IMihhHq9OBKMmQ8ddrdBApy8o+t1UlneX
EfpP8/rpKqHIx/2ZU7vzx7kFLLTnsjlpUYkOrToVURTS2pz2HBpLbvUJ0LovRBCU
1alNytw9GN7ZEPZYQcdODDqTDymLTz902+LgmRxtnBWYAFYvKZb+fCrctXY0GLg4
hxO/rbgGtzNxIATw8Ddo13J24tRKGCj8nWtO9q9HLqQ4R0rodf1oMUrRqrPs/7wG
mQEvaGKzJ4uAmesDbHE5g22aSMbuk5dj17BlKwku7XWVk5FYKlObBkd8vvqaLN0f
tfvunGWY38S+rp4MOqDKERPVt45gYKzBanVn9yQ2tvPI06A3qROd03dKwqp9UoYk
5vu5vbRQl+0pItKiy7IoOqiKwUOmLDNT5tV410pCk6V2mEXrc3A6UkvjUAS5c6R0
Yw8EOMVqfS95wyeLh7M0qXW+gSr/VYQEUDc/GSMKPxGnKnZrayR48lDVmW7loAO1
eL1OlPiynXRjTjFWul54BxrhI5sXGjryctWn2ceBzN/FI08qRYyOyTagQI5+n2FO
+RWPahCx5Ry8WyROLZ4z0jAbCEbyNJILilOyHAKAqCSO01dFL5jMtOYxyh9X4QfK
CYLxQ2iw9NFmfYLCVvmuE6MCUc/ktpjWIVv2TYMWMK4F3eEb2NwC1rraj0VhjPTt
WiIwVj3/nq7/CyD1hK/7NR/Ma/XKVbVQb3Akd56vXmntR4dnOIHEXicasyqozIMC
oOaSx4smEaDbKp3mvpiYRcaIsAN9npQ8gVQt/9XmgfJX5ISJywGpS+y/b36Vb+KV
IgnkzJFWjl4sE8b376HrsGbiyo811Vmm6Fn0RjERVw2ptcDLcnTBETx8E0dzXmHF
hzu339VPi0s78nO+rbdov5Tq34L76guTlqC/u9h9x2OfL/kjivQ4Lj9moz2Axu0o
6NDoqIyk4tDtjub7dvAhP8d6PKxAelLPProIjfYL7FPotgRa8dCOhe0iCHCn0ug0
P4px6o7bnHhDU9WJS1wnt9vx8uFzkxsQylewVFTPv1aAnkedpW8pybtNTUhh1cyc
ur5vNF5eabuObJ4v4a8bcSgpvu6M+8noUNJj1x9NyhiucJpIRcp6dPBmGJlnHaRP
ASzoTeMsc4UeyGdQRLjBzUTwj2cdznyoJoth5N1+l0c7tx+ffU6fuYnHmvWEsXbh
pAY8NNuiSYV9CaQrQQSPq/nqe+FWmxc7s6TIk1hJ4bsby7kvQ6/xM8UVZUb+mGli
1cyffCKKIU4KyBV4Ml49xKjLLNZ5AyXJi+SApnZszTIVwbMy+nWlpLjoN9airbNc
/DFryNzQ1/IUM5OT2mJkkEQNwkKOvNbnaeSTgpGkHqblAzifVDxYA5punKY6B/Mz
zMWAsfQi9nf9EIFeSptETXNkOBLOIATkq4Gc8BrPFQa1eIilMRaK6WENyFrRhVcd
6Vqh8vuOAG/T/S/LkBkah1hJ519UN6F1nVig6CNcjRg8Z5CxNfZR5Ov7h1izilNP
A/7UpyERlUbjO6ad0mRd1/TOzweS6VvuEIZTFl0aWlYHM421qwG+cfiOCuT/tQwS
xw1CcZkc84BKQ5kSX4FGZtPAHBcLoVW38jGbanRj74IyPAUXEwtzHlURM8QHgOyy
PfgePKJHmGK6hvLyRN34tYweyziaTQGBKWU4qZPy2v3ZLRhX/5xicG7m9Kq/yRlD
cRQpYdtBoLvYY2mteJfKg4oiTJCELWIrTtN+lWUvF/wfIe+U9bxWAHHmoVPMzHXL
MWmDk1JS1U6/lmOZaypJcaGiIE65ltz1t1aGU1m1ZixDne4BFsFndgKraLTGbbQU
j5n2r7FrWMRzFWn6P8NKHObhT5DFvEStlioDT/tLh3eRmz78OdyJTsJoHRAZIiCH
sZF5HwGKjqDE5KOsTcXc8YAp/AKjJMqXhpO1yHsf8J87w08wcbPKTU5W5Q6uWhk+
lHrZB3iP2gzymm+ZYmHNSh49TBl46Hwv6Xy89GlRjNwYNQfiREYcqQZWWK/kxgse
amIFkzQaW9M0yBo+o3rW5QlJihRU0BwKYouiCW2a+UhfLqhjM2r7r3cko4O2gPrt
pi9E0yogxxqc14Q/GhYrr10hpukUUyg++93LW+8dvOEQRvaA2d/RyeZRmxPfHpgj
PaJa4NEqIH9Q5EM7yc43+XsW3mEqANFlmXpxkjFnMB2E00r3l1L+oUGChRsVQG1D
HCJrvIOMb4JLV+aesrWiFsKwGg4CV3HfNYNIMbYs+KAD4zfG6dH3CKe31slhZYPs
GrZTTHlQ4vO8wLmph3T0uQRrpRs47CUjEvlgl8INvDh79Ttr9tExWOsjXeTNoYq1
ka1n2LbLxD921m1Iiwx0yw7kPOW0kXb7g0IRsqkMWyEzGNHYQy/9BL+86cODRCCf
POJxNMj7WOg6wqQShPnw3YkDOnsvc+WLJojDPOV5OJgWVRS5V8wQLaLh0aee4uqs
QYM7S9gDy5MQDvIK5YTe2iIJyehZylzZ1Hh+yoGqqnlwGCtJfpsW0iXmbtaqbIS2
o849jAmpXSQkA49LByUumaKl87YPKjD+D58uVfHQg/gDmqy1Rlr5uo2ZGqMdhxtB
MJAn7T0dUa8GmRIk8wjtJgEJ0/XOeFFAI2a6k1ZPLBhcPwh/TcFbZr3IS1w7B4x2
yhieXyHi5rn+zg1823jU8YUUHUptzriOf7vMPYseWU69DxAa9zyv8XaWkwiNDOnj
cVlgd01akr0aT2rcHSuR0prU//BoVIrlReRMjBfQNy/LJnQOlHt8Wde1mB2QDdcF
wSLwiB28AYnJEY7KyB17JWBFR9im7o5pvNtJCorEAH96Z9V0kPHAMZ9E1ccYvSHZ
6OdTJASsNfIf7PuGnZcLZsSxznIFuglKyi6S+MjONtDevUqwvN9GhssU683lA7FV
ASIau8f2jOUFkjtbN19wlz39AkPqW7e8u/mzdVHMd8NEyNqoUEEOQnmIAdhKUYIg
1ZMX4g/0jk/G9FNAITW/sLbV1ecQjumi6zjm4Fnwri3TlBNoGIbE4ErLiGLckiRs
dZaZxMn/kOkUXCVnt6KYDA0VkuOodWPI9XfavmfyXLF0wmj89M5JRtTVxJtBelx7
Qh+/KysL3+Waa+oXGsmcq2QlQt3f/Y3qrAthjUYOAjagHsaGOzjt4IrsqJH1+s/8
QshjBjAFbcLLEMbf8W0zFxghgds1PFTbyPq0n09g1DtKf0R1aALEHtslbhS78Fbt
kNhR43LKtu6v3v1/WdoIibzGh40afoPQXu+4N0BdEcaqdPqsqq7d+0H9oaA58EnB
f+9GH5PgItZNUH5dRJ2b2NwMMotnAqH8cJEzNsr6GdJT17b8Z1wX9GCYT970Lf7J
uQ8jkC2re1M85UIB/Q9/Gtt4dj6pH7xwIcR34aSX/jkDUp9OEVWS09Jskhb8ST2Z
50hlREydIRH6PZ+S74xZEJzBET4kXppBTcc4LtPE8PXWK/ikZYDRPTdJ6soC7YGE
/lk8uHXfeDsVhsSD1GFmAM+3OIiMLYO3VkFy7ze+kZRjnVBFTJefwSeKpWsD/3Ka
4kRAorMLZgPJX0DTmxCl+0Va6hN6rX88IGATqrlIZdRhxTSCbpDZSun4u10OLaJV
WcDAbttAnuvxtken2E/AN2ZVm80Ku7eswZcpVjOy+0QnEi4/obzgNPM0TfYf1F0D
bM9SHdaDnh+6J0ujmbSH1kNFk84vKUZ0VCvbK5QA71niO+ovRt1FWQKLr224mUlc
VK+E7QOWKwx+DzJUMouLkkIkCxrJTdR0PEZfhCnHYoG/lH6WyXBy6jnQvjXf18gT
Iir9rH5KnShngUdxx4HIH9niUEH1UJ7+c8XcC/ChziqySpvbVLHvnSCQxJ6vvJrJ
7lprAG+zEnJDIzvU2tHZk27GlIDdwAB9hEsrVW6l0D0T/Y+ONntdA7AJ8OP/Qfgr
O2VG7jwRwXgdxBMfTxRz3F89asJGowzL0bNPj8sjDVpW1P0shOJsPClOPHbMOdz6
UmNC8dfE+O4hoaSBPDRQSyYHnbre0rl9ND7CGl2oqU0aF+3UJjpS1PPUTFJ3eX+Y
118/bIAeVdtjsD3pQ+JodDj13QIskDMX+cfPo48WXz0YCJEBkqQOcRe08akhTR8q
uW/DfF/sSO2MCeIKpquDaOXpK52vxB27dxyr2UifPiSFlzyTLs6gG13WyHVJybmI
1ayeX1AVbk+7xiCSlRMBFxOEYNUSLgpBXihavMxEkFMDE3ZuXmMKOEwZXBqOHM2t
FQxvuD/V2mTHr6gzWM49h2udLZL+lofzo3MrmHu2FIQOP4U614sOm1S556x/rLZa
YsR/a2LlFbMMiWu5z+bq0WbmwQ89hd22S5RILZiGHOZkLsbiICLfTngFvzzrQGML
Y74F+uGOo6a6YzeI38hEPxYb1itdVCOvFBRjybXjVuYGzT+3zHmN7aaymW8wGbfP
eQfOGBX+VLfpcHJqH+/NRWMAOaCbJC5i5JMwgrI8TqEDCpTmFk0zgyUQcjbDpVEU
VNfW413Pfepc0V0U/3vCInt0inHHr8dGkQbi7h+sV3ydfBqrQE7W6WfsAM5y25eP
Y3a0WjNx9IyfR1ONWTQgvSOySabsNu4eZwsWCtkS61YKpPUAfZr3ip7BAwy3tYau
JEl3EnD1OkIxPLcnyeZO0zG6tA7w1uVyJV2XzpaB3oIkAwfutHAgJUjMNWF8SCS/
bF6N+C0hRZPkRBEjjwuF/0Iz7PnNA7fI8mkk6B9d9rIDfSNhABd/5HOnf6t8fH87
4Oh/fpIrva/7to5LnVWJ2p4QiyRXt6nxUHhNABNT6UnaMpH75cM6fiu8C1q0/zBc
EutFmKFDUNUxZHxUU71y7GkaAyd4BnGG8jaRhldNPdBEnN8JWHTVbd1kA1M4s3Xo
ICdJsKtDrIcDhatoUxE1Cx4kY6QNoBJ+DHgYjvPek9ACYQDDXXjlNnUA61Ev7w+S
Sh5aOwfQHRAQvAUh0Iqf1wJ0TTG74xsNbvJIJlqzfViPwW10HKM5h1+Oa0evOk0l
ZeSS1jOaqZGT4K7SPqa6p4SdCxrsoiW5jC6IBRBi3fj2yg67Ln+ZExMC+FRrVV51
jm8/fI1aHVQWGtKLDqYi0s5GbGRqRUFg+ttHJEqME6Su7+59SZTdkLkS250O1irP
ibFTHOB8GDlti94+xJqUaByC6+vpjy0SEECHnNoksAdHMKnNWB8hLhigItq+CGlw
CYl3lsq7LiN5ynbEHdhrs2/L1d/lfCxQT3cXsqjf/REK83yBrgwuGC+ge1KY6rhU
o60Sd0ZqY63m9c+x6IiwS/hqhZBc5CL5cJxDH80dwqU2mMYd7DG8Qn1zlDykDVc4
ki/kXp36y5QVoBEXEqfRdaKp6npf2HA1A4xyB3vQPbEp/AFgaaWHQ+oiYkaelaL/
AsFJUb0Tou+vqA9c9JkhX8I/gTFCsu8NPIqYVdjIKWyfSUpToc1o3bAfimrgVlpD
rhgKMAEPrbPVRGm1ziAsn9qGBngNtRbwjM0g1di/ZKR1KMhPZERkOhgJl1yLlOqC
p1ZfzjwhzkWSnzL0gESXUXLEehd+psCRHbn9CLeNKXBpEVd50AMJUFgo2W2Fsajn
xTMPMdmO/mHiNSD2deB7mM5vZhPNENdtaCZghLljdbSDks3158VoBpMDU2X98QPw
2Tqa2WcvkLbCJFRhfvISfzEf7o/0i5NyR+xt5XYe4y7LR/gjbdKoaYDZMWkMeAgR
TDdTgexULu42UcbbUqfCupjsisTrbGEMXLZ0DftqtBV0OdYXEIbo9MSnSMxxBoXX
EcvoaPeac8dwEqDsNeBoG2l4EiCN7MQ9T/0OnUKsfTkNOnAXMbpFZXgToJTCOJzB
DfYCsbBGl7WFc3OsGd9AkNzAK6tRfL2Xc/e4e5JYvpHFR8UjLcNq478koreQ8k0O
QPeKHfYVwbqnU/EIQYGzHC2OG+c4Q5xdCacQ+/r+5LQ1zSAqDCkB7A87HaZhcagQ
S903vZiXYL49djPzxU9OawRYzfzcxOiWpIKxKzt4qiC9XDarRHWNSMM1Gm1hGFx2
rob3PRfYNkV5VOnS9yXGvatkMwGS5N07n/2Y1oifNnKADKdtfZvKJfTXsrPZKjcB
R/MNUrq0dlWx/DTUGVKis1lZtoX1YUmlC9OyFvowntU5VSzZhUkgrONc45eUCUsq
JGFDxBIK9KvDKdF56HQb88wzXqrA/x7/QDGBcd9hsPgjiZqmwtHhQSFIksHi3HyU
9gixYXxI3L5GqILzrrvO93oZ1l9pfj2Rc4dI5I4CQzm/o1jx8NVNi05+gykimcIx
dKM/7k++sb3vKI7QAy/rYJt4wXvHTfGbPB65OxRHomKD2WFPXhzda9gLnKf/Gjix
aPEK4optZ7kwfndqOKZJifNKJ8qW0XjYxDhd2lUJPg1a4cDSbgPZwcKGk0J8DSlq
ooE5wNA5hkwIP36y8JEoopcyBXe/kYJpl/7shMq+6b+J9M6VA4EKceyEK8vNu12/
g8kVZ6YywNj3O4NookoI6IdealhgfE6gpMpoZ2GKIhLXTjXPFGDQSP5qJ/fidVkk
LIeghKSe5IMx3/UQncEX4OLaPdC5hq+tUCrKXTlkZrGGAOi56L4AfHjmvinG3JKl
yT726syiWFo0FFVr/DrHlOyYR7KgwLjP1M0k6+mkArh+4rOG3lLiuSZiWE0Zb+xV
0fy1tG5hfT2AEjLFB8vnhbcY/8GyR632Keknil21wQA/JejM3p2s5KTCTcRQ0/Zl
9gO4yDmNzaPPKRJ59YlQ0lNg+YNq2X5ERHgREAX/+IjcOE8HmO9EIJ8Ngmlqtb/G
798cm/6IXqvqsaDoUYxDaTwe5Czxg8ej8mPPTewobzc0xdRd6Y8gL3lz+XZR0IK0
zQLjyawt10uEf1Malq2SrX2zZhlxwMVQlMb994daRJqG+aKthba9V+aLVJdour4I
1vUA9MkZzTnE/DdroxPQV57426wjVv3Q1txHC5UcTfa4d4KS+khBu1tZ6HqnpCqD
XaH47cI8qmC4UIJn+HemwDnygxTU3nk7KtNe7QjQuN4HnCWGB6MRLZ9+Q9m0/HOE
oZ7v8fz5hGiDtQ2dbyPdkUFRXM94fXww3LX54a6VEsMXlJ8WJzQONL67MWNjEw1z
4Cy7kefZ8jPYIHyrcwZN7d6xHhYNg7McLpoFa8b/0oS/eiuv4MEiUj9rP8FcsKEJ
F/Vkxvge73AI+pcbh8EL7GYFitGLUFYigN6BHt2WoaLnNv/sAL1Wj1XmOzM90Ne1
eGuBI6J8x8VRXRLxE3YJ0A4dfeQ3/sRqv/AJIMQkM+btdaWosUpLmrLzwDBar9KP
V63K+hGIOBchI+X5IisNVR5EaVm6zhNzREoZgSTR+3xAXnHi3MhgRdJtkt45Jxc9
qMqIb+wQxQmawukIon1q4+xrmyBImdrGjNIAbsS2yFvQjASNPQyG+dWi7TPv+1S0
iJXo+ayw6Mn/QNhNmR9Jl5y8RxTdGao7cv5onCQQUQKEQr2+8H/UE14wMOrYpIMu
sHfef6J78nHhA/uHpiUONOlNH6WjN0bZe3FftvELlP85q1cD6BTeWbsz8PRxxDLX
5rIc2c7P4a5pZGOUu9LwBo6kByKvS0LndfT8OvQEmfr/x0YhP5U52SbRgi5/bpt6
7PxqZHtgh4jcJbjtARU7jWuZ8/270LVLHTDQU/qcHEMEcS5gMU1WmgxQ/bEe+xRo
572cmVCDyC0bYy5VkRgX+Rl9gt6QTscL36LgZprNaD1s1HV4aVf5dyIoF0aiW+cT
OotY6dmfrPR9MIdt6AHVG0rX5NCdqIsUfwV04eJZh7cevUwVeKeADpNP0pMoZaxw
bdEq+Sf2BE/O5L2mW0uHfRvS3CBw0LqM1nwh4mBymhB6xtGdN7DAZZAoPdKIW97W
xZsUwiqnJkknHzzElBoai5iLGoTqNH7QNFilC6wbiztf4XPGBJ6jZj9+5pJjp6qO
04Kz94nEqvudq74zviylJyPjOm6VJzBhbXasuusJalovqpKRDuJdALqsEd693dwj
JbM8hBHLWT6lJ7OygQRvC8sjr5f35OnvqKdMcSCPj8L0VbTb7o6eyE2QHbBcl0xt
Kl1NIrsqip9sQ6jfOZnD8kLMvli+pHPPoaIjfMWPRMcagEAbuTb5PjqdWFwpnlK8
e4oowGu43hHviuK5ZThknKbKh825AFQoB1BoQ7HcwFyk8yJ3PgpHE2gRT2hRe+D1
kZ23mFAgNuXW4YpoYPEwA1K/VWOinos4n0IMaaFuKJl+eBMvU6Kw8xNMC6OzPlso
MsBYHu01tE3B9RL+Zu4BJa0wM/vnBA1pXXHUkgrjj17aKluSqlmGihSSpB39LBTr
h/JOhV48shHzRjrr8NtUbS3AufyoGVu6lDlssg78V68adrK5vYyTsxZjblLedf4l
On28UW4S8KFOR6UyOrJ4dIJNgF2b9Eggqm9NPM6EoV5NM4Iwu9YtJAbTelScqqDB
ONLRma9daJSV8WIpgUT++f0o6MzoOPr5d40Y+UDFjc06vNLH6KRxjfLIw7/Xh85s
+pMU6gxiqZ7afwf2DQdXNPyJ9k1s4M6dJYrEAOEZaLMIB4oT+P3FUGUnGQOBCwmT
Wvf43VnJdy+Yk2Rh443YiF4wHLVvos3LKW8bbS2RYj1XMwaZW4huJYRB3KicU4lW
5id4WGQEhvYgki1y3mlimuJHu7DxCReb+EKF0hrZ5mKLkSauZsaD2gGgZU+ZLKzo
zX+SQJ2PbFRrBmJCjl6RQhRJpibuVAK+Ei4DnU/pWaa37GdAjYaaqieszHYXdWZZ
i+Z+7AwxegOrZu959Czy6dt4gJPICXHAf4yef/lXpcv5lW2Xe0IJTbpUU8cMhQkH
8RoRusF2XxwVrIUvjV+594mOg8dZKDMTOBSYtE4eM5QtvD1L98HUaKg+whGk/3G+
EoWwIXMSWxvnOBVbeydy3/z56Z6zVs7UZLZ176hwz9nbNnIAhaTWDzJthNrxWtbp
murqKesFs6kcv1Cwkyyzp3r5UbbzP4mD+q0Vvkd4qSPbVhtPILDkuqBoH9cIH5Lh
dimhTBpgRQgOIoXW7hvLU9ogH/JWJHsQsc/qHRcek6nSv0pCTE524cpPfMdms4FE
XGGkhw0F9bxU6et46hLSaoV4ApREqPanGWTBUEWVvol5/WSUj52E9sRU4KtABLZ1
GRxfyhXu0T4YNQc/Hw4gM3Tdj2QfcEtmdQWTgbGohCLvQJ3kdl3YyhJ4T36J3BKM
BpprXYp6ub7tWBms0LTRyJuYCBCwzDHWFCucOdNdoUkemL2UaGMrhIBvKGDKnF6r
c09YB9Q7KT8rG+U655KVw+lD++A/MSR5bbc6bQ1+Qbiz7w79FvGPDPM9vPFb6WGl
z1aOnHYp42PHfwVNyWipCBC9foQwT1ZvNtXK0YM/KpFWAqfYodaIMiSpE4X7GsvS
uXitz5kp7n+DPkGtgcoM4wDeFR1q7My3R0eYuSKdow1QA6W1Rk+gARTAztMZ8euT
fy0zB8jY9l8p1e6DsYSaGPMvoPdWYkQWxvkfg/i3IdvWkNCdzYTwFReprczKgxh4
P8oVG4meQMAacxtxBmKAm4nhsx6fFtqyLAqRUVqSlVg4Z6fE5XB5vQ2f0hnpSzs/
lrHUXCVCPhHTf7uzn1S9O4ypEsIVLcbsNdh3kh61zlrimEJW1uuqHJl5OYWXqjwt
BLGR8frr68Pfpbou3VFPSmywvRpVR/hA4gXp7cWdSwvcDsmUVyoQSm8fAeBeYeLW
qgk4TkrHSxv7T2Kc67gtvuLWY9yRKYjwN9shlaxtST5YnT41yfVsx/m0Cj6ymJtU
nfdDiM1ecmRvc5zwpwxZR+RwvFEFRKBNmD2GaxevVAArKz+SSYyaLIWwMS0jKSAo
MPFMeFwiKeCLJ04S5H9ptC2VrWvH3zdGqXQ6q1P+XqL5TL50oMoPft4WmZ0+CvtV
wkZ2fqMJQ2N83XyVzmNN+/CTZCJx0GV8Kkcj66XLUSyLotBAFsnT38vTIa0iiMhq
RT8FhDaeVkJI+FX6bEOKxTYLPDL4QRzTgOchQJ2mz6oUMhOcp1ppQqD5vuSBrm04
nLtOXlA1joV28Wm2p2Tj/u5lEq/F7kyKRHH1kjCivysNNlOnb1lXrlmfbBxTg37Y
rQdP2Z1w8kES77SYbmD4iqfncRjuvMn9uZT0QXkzDgIK+3jUAMnyobPGVFpLbzb1
uDnlS9M+bK3SuzWjLOAHC6CMJoRAZDQ9uJZvyECSErQ6H5fwoEBIRSVcfFKTd/+2
FUW+CPD3Tx9YfDNTXHSv48GEFZnCnvGMVntuEcG2ihJA/4OKNRmOON4Vqd+gIskh
/UH4tJsvl0OHWZYtHgGK9wOkcCL1iB9A7VFwToNNId4+BxBkoezppgK0rGKpclCG
n62rX++34WDt8mN3La9Y9Gxsktbym8vaqqRcJQL05sm/Kbg8co9iMnWl5vZMArl7
Y+kXghNGukhjRZa5In4OMegg+Mx1svaToXo5uhFHc4EU7pOGpTuBDUmhqJkCK7JT
+4p7VWiYoh2CuF5WEE0qE1k8zwc1oP87fyuuGXkOIXpt1BVhtWjr/sPmGhrb/15A
qmw2oEe53prZhOh9Q/fIRM7I8giHiOQtC4v3t6zeZZjBctEmNduWPKt+yzmYdii3
n2YEy8xyfag8DYZiS8Pk7WsyN7Z0UjdrbRlVloVbUdAGakJ7S6YLf2cZSrapmxDc
hJPntzeoyyT7DpsHlK29wSGh9z8hsL//zchfa1fgK+BncGFI0Jq/1q1xNR66HtGR
N7gJVuYCusOi+kt/cQx+mMPyHj/apiSgF1xy0jepFL4vhixrkhTTD5eBlb/OdnIZ
AW6lTytMDhaUofvvBRtBl6pXNtwBT3IlIcxeZ94Y0E8Lh7p48EoWYsxY59yMroA6
9GzgnzRXjhn+kiTrrY5VMv39HYuvJeNmAdTWwlWH8TbwghV6d0K/Jg1nRDeEjm87
1qkVsN4xAJrPJcWAe6eeS6HqUNqZg+4Swpsaqc3VSOxXB0L+WGO9TCmdxdNibfBZ
6+m/l50B0wBAubIsJVm+YYqLkeyXwuZ+YS/E52qNuFDhb4yMqT3F8LUWUtfMMLB6
+r0VxQTjeJMP8lpQ+NweiIa1jXkXcKoxPb6Zm9uD9IAOUsLFNY7R+vDGSdC5E7eI
59E8zl5ueo2Qe0BjZ0+k/ubEGWcfbUt+h3gbE5KRSaHux8AKGlucEbyDe54S35sE
xSB2CCBGiX+kdDmYlyoJ4EMVGWW1clRJS70IK+HFywfv8bM5Q8Owf4GjgC3s6Qay
0RwFAmXOfObEHx/e5bYbaPSLfU5HNND7X0/VLfAkTS+QBxodTKlFft9wpHTty0zx
5A1rjGWAEz3nuxBx6BIq8LJO9LsnXQG2mp0uzxJN0zSrKjcznqDK//eps/Q7BscW
XQol0tEkVwvPhmlqG2/jwJqdk4mp9bOqIU62MF0Z6BvZrxsgcumEeRc/OL6qRMis
IUuYAdPFWLZWo7SHYCbKxFnnanTWxwvwq0ClsdFdz+fNS1zFwv06XRFYQuIcY88z
9lM45LJ65p2Mt4IHTJ50dnKjFw2VlhglTzovYnAC2S9jMqXHPRMLznE7o7KO21wO
LO/ZaHJHIwflqpLyesKS4oiucSu9dFFuPdwibbT0vlYK9aA3ZrZMdPJNL0u9RoZM
K6xdFpXVgSjwJKQ30vO1WzhaAJRQ8LOhG+jVqeTCJUucN1hLO3O9KrNHiyaxZbJT
2C5FZgk8N24x/wZGs+fpF/a9MlaLqEmOqLKPADzbySNInEHYT4L97UJ/ubPgpJz8
g8PGGeHBS2lfS33MUrDJAo4fkP58K9wbKAyMfamts9u5x5ADtAPNcJSxok2/3uMO
jsJhKk01MZsN7X9ca/YXtxcnxUSbyzbIgRRgzb3LZrkvW/OfqKyjC6sd4HmnEopU
CVPy0b/O7iXLyP8D2IY7N/P6drXEXjuYdHkGErDIKcTegVM87cEXFT2guKvoZ8kb
yvPadEBpX40u6kRdwGgjgL7prHEG1GUkCJICe/jn2qKmZ5MNrs2vS4dgswHQcKGe
7KT0J5uunaOaSoC4dKgAP/HfdcVBk01b8W8DWyYenFEvjX4xnNJ/sULCPuiPmjZo
xMQW/JyStG/Hz6882V23+ZE+sJF8f9Vl04N5OazuE/wd9vkFEHX13ii2h7cMo1hk
Idoh1cpbTUzqTxjUvQMLjw/Lz9vakxhqecbVHPl+2XjTTHz4beWlosW5JmC4Clg4
lddy0Ty2FwZ7qzfGQH7bhWBQ1A13Mipa7oF1RNkq1SWwABSKgRpLiy6xOT2haA6b
17SDiruGgeYWI35OLDoJ+lB7zQtMkhHQu92b9A7l4F3fd0lm081COuonwzXtlURW
c++TGMGmIo2+gxpoPMWzO2tWd4pJzPV5Xvh+Lz5ivx+vL0P6ftiOKvs2SU4wwzBw
jUY8rWo3YiLAGhthXRhoNY7zr79v1mKg5JE4i5J3rn1OKWWx3wnCjqZeCkn8SqCY
1r/v+O8AnKvWDsDQgnzbDWJNrXAA5eF3XzqIrT0DpRo0z5BgsQ2m8okfc407trJa
IRp3BwHH3ln+PNXCPgBo3b/NLz9zHW+1EpomNRMzBtGzLMXnAA1WQT8Xh1P8GlOP
ZluCwrPERW2S8iv7UjcTujONyfZIDQGlBolNL9KiOXKzfU9GOUZb95jwG9IfQcu1
pbXE7vC3YNyPktJOtWHbABrjBOv+2wAsDXW4An16TJYGczKt9ss1gXfeGUI2q66d
vNYg+bZrS/t/FZuLRPAOjYXmGCjxKPMdbK8QhDk3Gq9zz2m+nhzJvhUxhIqsdN1J
gQSHgy/g5mKyxV/TFVgZP8gWQBVc57OKhz5vyQMJhEsOMw1YV0BHAFcyXMstq1Z8
jBGG8rw4Z1JWpzf03NqvGX4NyKE1vm18PHrytghS1YZTgROkbrmDylJoebHz+2BS
FbnMJu8oxE3TwhJbbufx2yH20sRVfJ6z0yj1Vr4B0S55xMUwajU6QHEjui52YyCC
0I9QPVtvoVO8Q+yA4Rx5OPQVSfeX09etfDGi4aoTP0gdvbpS8yuigcMYnicPgmdN
58IqWTfWOHq7wJ7gTa9CtQmQMLu5zmSDp391C7p1wOzCa094zZyWsblDvdcXZJy6
x9Xun+GSG14/ZfNV1vLBglu2gM7Ni950cViGnMPG0ILlf5MGcj7vBthzg2RvOgg9
f/R+Goo8ReRBYDmI4rsnrm+8ncwo8YWnpPGhWa5L3L6DANgLeMwHE735PhM8/8oE
qFBWPzW9ldMjxm4ernyB4C9/ikNh8N8txv6TinSU4SEieA0wQi6zzfPN5R5ijWAQ
J6vSQdYXq3jSCZvGfNQvIIaONnRCagKYnDZzXQGjRaeNccV8SWt4f7JBWo7sGjsF
DhBXJgt2Ktre41+S+lkscKy68aElsiMtjKh1hXwfluBdKyoEdwvsmCq9/OHkBVMu
Tos4MOvOLZZj1aLaBqmt1xaEui1atM8n/mH5HmYcOZWqCJBtVJDZgrUcKK2X3C+G
N0rMbPRWlLm4R8c5Sw5zDbrz+RwEEsBvVbF2qmKIvZDxLKuPlAXOk6TIOSMn0XI/
4g/mxFBJPQDFZZXqferu18UYhRUU0gyvDWcbfYToPWjztMSWNtExn7DBMKEGILOc
yFiXUFqk9Hmw4W6kkNdZLXtKL0WArHamGxg5swd2XVlaeYOnWUJUb987PSQkKalP
PJFf+RHMvz0MdzS2SZLOm4VCVgO6MLhG0ybDwGFrAyhXE/tDNRQuKkZ3LlQ6+Dgr
S0EHkVECL8tApe3y3z1E1td1fuxRK5SaU96vJJCaZDnF7zQJoNyRVABop2YdgOrq
4VrJ+bIkN0R5mx7wddbu2Cli34nUazumZ9CLN6oM2PohrdYKR5p0oCMKXYV9Eko/
iu1yn2lF6/sEM7ODyjZPFjZ26bKZY1SwQK6uFRNbmlT5Rsi/Et9nc3qvRmWSLLkC
10GIAbtifGZpPpSsB2hc9aqC+q1hRPMB/bV0Upi2WpzURO2mGTQibjq//Lw/6W51
6E2emxCRy7MON4FyQOA14XS7lBwvu8A1frohitPvwD4kepIbcs2QcPmKgNjWQh9G
ShlOhU+Sa8ZYAqRKEDvOBd4kKIrQcOIsnuBrLA1ltkR0fX1H/pFNXDw4kqB5T9+D
DDbgJW86kuKNA10zK3BIO3pq+9KaA/1UyQ7yVLzDD01jS9hrmSB6xJZDbYpHxn4n
+fwJQxTsDfz+PNZFt3RMjzm/a0orunrL2vCaD3W2wvfOOgNRxsoM9Z6l4GwnpYHC
SGUBJqHsBM+kecfvWRAKU67Von5cKfzzYQx+P4ADM7/L+gf639Zg/aKD/6IweKyb
EwYuyB+6pPS4I7NQHTYNqF1DTXA6m64vqHzIUS9dRDFP3admNGkwQpq1IXAgbVts
r9wF/dRvy22pajBnjd8hU2qMMu1rDFKawlOXHuTOq3Q3YAdJYS4UvDjJnnzYOrs4
xdqdyT63qsy6Sn4fDmWSzxJeYyoRlSDS1unqa5WsqbJ7V6v51L6QlFP7QNEI3Fv1
FN4txWMZelmCrtACUPsUDwHtLRUGqhLOKwqMxQ+3pH3zoRjzdxZLrWyH1g8Sv4a1
bIS03SZUM8xZ3tFm02scLt5ii2JcXyq8kPEqZc/K8OZni2HiGdx1BQTwoc9McHCh
gjsUJtF+/9fIs7aDm3Yp2aP+h6YvcdQJLYmOYn17oUbdzeMw6+ImjTYMLBANOOk3
TrhxQ+mzOXb0Z24ih5M5GeUWpjhdSuf9rB0kztR+O1YREDxFaOkFLPkoEknTaoHb
znC+2pgg4U6Xu/dmhXnLvgs8azk13Mznh+aLtiLDnlcA76OGADucDffLWB43myhr
4GHd3loA2dNUaX+9mQiiOLL+uQDXJMvJ/Eie22r1jcbJjXZ9pQPh0SnjGkaFXfqn
IvJGKkngihrSNOxwugPQMexBIi3TSIzI80ZHfxO+Y+DFitepE8rCS2JDukFR2cIV
RRRt5GtOy7zCcDNe/DRrfPB026dJ5uY9/g8SnZ+hpQkdY7AHo1lTQmXFMFoGC86M
baFWdrFh1i2BBGkOFDNPzi+W5Uxx2ijJ4hSIS7fLcUAmZLiujLrZ35lv6noN7XNe
cj7pA84+o96VZCy9E4yUgZK0Z+rpzoB3Cen5wppEnW3rBYSGuX5miruqbUqgW3Kg
XXy7fpQ5F66ks1MIJxES0Fo0sCFivQw1KC4nCGWNvpkhMmFeRSStMw/+PbAfqdRb
qg9jlp7e5aO6M4C0JV27++rkxCTT0ns9G1lx2su4JpPMfgA92JxLzMmNcIGxZqyt
sHo48FW50PJrSa4lseektrG0QmjrdDNYOU46pVpkgEdXRYJpW5KMuyG8d/h7M74C
L3ay3ykbmU7M0jgmV5DiQpah74hd86W3jxMJ7CoaFD1UOSSKcHsdMak2vicL5xGN
REXWW1AGSE5X91Ymb/CPKmPyJzSQjb8qQ3LyFX/X8Obuv8wyTstmnpU1eeqyWRl3
5dC3IgR2UltvUUlP38T1PPrK1XfTALEj0Q/QXLAP05GF8m+g8TL/m6UtT/KZLi8T
t9byVAWb7ZnX0hlD9rduBVzsnAVqbLTME5+dmt65jE8TI7juPnnbDMT4g+gHhl2r
QT5VhUUXnOu8T2qRbiR83pMC0tjoaulQaHWC9jL974/wnoCyjXE6DdWZEMrLMs63
DOZElzCyGMAYZI7OgBQ+RoXk5cH8m2XnCmiCQssmTq/+ZPJMmgBCx/yw++PtMtzP
u2M+UjTFdcues3WyPjSB1jaTUcQGVm103xzQzY4u7PeLpCpyoukYzknzlVOaOC5N
+uauYMBW+kKDy8ZWm/6fUD8wb2HFfjwzygEV8iaqhQplFy/31PhtzJzI+VavabSQ
YVEjiKvNe8CwPZn6ArCqnz4eE7R6Ibt0kuJ+JWeXiG+TZzKMgj8b/GN6w1hsj1er
/ya89+qJfKAjFKm1XHaV91usdhiP9IqH/Mxp1+FtSBjTqycG4HxlVy/MjLHlOL7h
WCFMPjwI5Z1zYumn2qT9pSlaCwik/Xn03FFU1fOGr0/oveaEKFHgWhvegF4knwSx
CwVEqNK4YxvtQXmieNZvxcG2olzDPqFGMWP4t+edgesEOCf2QVmrGFgZ9XOub1rG
rWV/unqZRwOd1IbN1nsRNZkFTwz/nPXI3VqnaUO/cv7cTpuKdUDj7UBenNBkTGo8
xWX0Dpx9I7Xrg4lZkwB7rNcB46qyS79fqAbyxAGM3XBG7jLh0quTufqNsRVuAjvU
g1MA4k3T65KZSvKo47eiY9nnTMKq119AhSr6Cfl1BsRSeMTlCAXCATJ0anx9hy96
Plfm50a5JP4Q6Mu0HzW9sU4tGxsYB22o66oTN5/9Kpze/IAGZ/hJSEuEm8ABVw2Z
DlKg43XL8i+89Ol9oEgHWX63Q2T3wMOelcQR2/J2pz2kJcM+5KP7O4n31+h3UIdP
3sKdm9SoxqdgWrsEIbov+2sY80AYvUPnr8rCfpmErCjBj2guXRCLKSW2MRX0UWVn
z1psFrfmx9z2C0nO6MYYGYJLX/dAtPMJGtBP5BXPUKNWuEp6G6NMZX7t8F04rQBV
nKebiZWN7ywmDaL3NB3izeg1UDq9UiGpEWKQ257d3P+MQo3d5W4v4sTHRa5rVZZ9
akjJqD4Tql/azfmd/Di68Zv8UENeOX3vmgQ5nGLxu7UWRwbUk4PYTsovDQPeUMet
qn8iPUeblpalzetfmwRdiD5zLOUUtUjacD86TGmhOiwtv4rXSSITj1bLG87TRXmU
0TD8phG2SMbW0Y9pkePSszp0f4VSzlQTx862+nx8MePXubiDMaAkpB2edvLrTd5+
VRWbV6E2BBAn0FMVVX5OWFjFGZsuHgU2mzl8OMDXxoVNTF60h7qrUtABUjA67kCz
zajhpVfAdL5KFSX2euc9OGkxJHGX5dEMNkVD/bwMnmC6GkfvBimdzucp1vB7wy4M
wS+ZVfoD2fl/Sr4k6nYf3tK2/7ZKQPWGvJ10veG2ZFDyGglnKSzJomLTLdNi256s
2pEr2u8Bwp+1wDFDu/lCH/SR3rwEEe+cNbEUUpXF3GGA+fXQz6vzPS4v7nHfNt5B
wBTtj4zMHGwNfpAGqcAidZHaVmWxTPWgsKB2kVHcEHq6HluROP/frKyYX1rtnIM0
OtztRCLJibrMHqAZO131Jm3ADah8ZVXOQTGkuxfqHPls168uUC0z04GtxnIuTsso
0tT/BkR3jcPLjlRyhpe1si3ZJ3A4qrUzC0vMNe8s+pdD5HLelpMBAk1VW2EIRZ+D
goJZoJtLZhpaatS5P+ufSfnHeFfYXhfF7WMqn2zrq9WYUKP3ZySaCr7eY8OsrwA+
lAJEnTiVtY1FLrciyCLudKIhtj41zebH+C1ERyjkYJqRClejtRuJVwLxrayCfmKz
2kb/zB9d9E2wiC8KqZ9apbjAFJUIcsTnUQ9QnSC52RIS7Ktzoe9XbWCYUF6M8i0N
kDMaMDXWtdeyedZ1wQ0iT7jAD9jmJGPPXsGBfWaAO+CGTmKPf68qsYCQBcjhoYPH
pbWGdfbIdXmsLnhWUm9jZlKhGVe0PD20GPT3Ssg1Pu6Qe4PB9NdMONTaum/FjIyo
pmk3iKbi4BlVNxRBfLeO0GFZzKuKDFE0oCqnMA+6nA46q9kypAvyElZprA8olUd7
3X3iCQ4GwevA23+bljez89blSIeMlnLZLe+9sRQSbfoYF9RoLjZY0mc6y2jDdBEH
d7CZ27wjHPm+xsvJbYrJsTzQc9tdET/LrommTF3/17tK8Q8zvcAgCt3FSjR8DFGO
GozTQ2AW19LjNFTgIJyturp8TotEjU722dDhkpwaQCndm6sDlK7/sIrB75a2CYkC
nI0v0o/XjkxbPl+RmBIkCs5WLT7V9Z0kiEvHUTqN7sHSwPfFH6aHgatLZgdk4vtm
Y5mSaEfpfdo67D2iUNIKGmmJc9kYYtvi9kRw06sEUnfpOkgbUyM0HPJnsfYN22Dj
zxDhaUg0cO+fePf7okSBJwtWJsY4uS+5IBF1+AGBvfyAUKs76L9GoLN/39siDgWz
LLOtX2qAHRh+Ty830VBa84N/TZ95WQSRVOgIfpf7bBfL0YbWsnZFQIFoDtGHr99/
rX/tR4cpzkWhrEpEe4VAmj1BzrDAlJAQNvb0iYYFtW/7K7bwPbC/f12YgRDsYRrL
nQBQkbNQmWs339Xmih9gkpQSivz1RxiWTP9ezqOvjIIgK70itscv3wJ7FZK7QgXc
nGqvs81wYGkaLY2cOaYk+W9FbCYslTEkTn5WvE5v3ePxhbcrWe4p4OOnJB19iPje
WjeOdRoyX7lnUhAUslWWe1A/I6YVsQ4mXEyBhM9oUvD7+twgkWAvefm+75P9hl7K
i9B2do/3FfEldtNnvICojWDNv/uB5dTFhAI2rxJVC7UubWNdMY4kjJAtKiyk4zTp
lw5xiz1MuXpPLea9+fHDLmJEpDCm5xCRCO+ZqMhOfH7ZsDcMb0xLjOyFfSpwlX0U
iV/sClNtfNOD5siAyS+l5vRxLpQGLuo2SpxeiwM6iaAIeEMhAZnZqDoxzrI7CBLQ
+exKI4pQQEHxizcLRiAy14jo2hr6B3UBl1Fc/Qr/zkyTqu3D57xXD33tlXbd9pSo
Pk+VT5YvcZQSR2xjxgPywZpxZEndtUiUXV/m0XoJQ1QSPIouOC8mdaaAYkA71EWE
fi+pE9KYALUqUMCNwggXxmEpPR0+wS1N3ukE3AhhiTmbPsQFgaqCzCnG9tRwd7Xx
Gm8gPRpso5809sk9xCvv2u1e15rn8fQU3Mt/y4xcoieJ729BvmhSvQGvyYt7yB7/
9bUoEJ3U7bVOxZ3q0jxe40mhrq+Q0ENAdbqk8ekhdqVfBCxZpO3LOo7tr7O+8Ykr
iHov4E6smb9KlEnFajfE3255SyWvQnbqv9ocYBex3M5zQ9qMKSVt0v7HkNKCVMUv
fvOY5hwc8moJzllf1flgUmgHuE+4+082BIIchm0Qu0QVUb34IfDqIbV+U0Ardyt1
B5mN+LCQg+yUfvPOAjNZ4WxY9/rSk73lEVze8OzYYpoZ8PVh1zqr4rWR5nb4C6Wz
OJ2NNwjDJiUXddS7h7lJ/Wkm2PhWrLFA4MbrWnfkk/+fNBXD5rWXIycD4k9DSYQ8
33XLk9H6EjiDUIwA6dBKKRJbOCkAdxUj3zPsqUL4dQuAgstIWVo8AtxmBocJ544y
BvKK5rmj3HoAnLHz/arpUGm0+JZLdllc04btWxuaR6U9IYtRSP3Nou6zj/gij3DH
AtSvo3ZY228ReufLi/M8wSn9okMGkQ5QrVUF9YZ2BHhqJ4jQgM/YONK8DgdLN3Ah
/vZZ5RJ0eoOyj8esABRZdyY+empbhIhKYKT4/88mG6Vh025lUdUQjRGvvAMHhLJV
aRwqzyPLAtbcJPPmfzBcYv7Z0NEM/1ZnHA7aDcooMdXIBCJ8CTAkyIztulnAwghG
r2LcevF7UUXZHGizoNqN+r49bYReLm00OYt6tfXWygJPfnvNAZMiXtIaXu/NbqmG
lgdS6RjE2VdzsGfD48/EMtgu5LdvEj7Vb62UQHRWsXQYzpq7pJ7EKNvTv4krS2GJ
Eijk0OA6J3jdk/H6c7QqBIeAw9YWiRDLodtEff6sqN9UH+gByI+BIhZtUMIW0Q0q
cGmWuNeNv6kb4prEVn1+FKk3qx21kln1W4YQkgUWWhIJzrqNqX9Z2TaxlEi676ct
RZvYebO70ffCeTAm8r2RNRvcfEX/EUypgGfk5I6tM7rhTbkclbiKWL1Z06l/E9/z
JtSmAb3nsyOLQ0cj2Bfaxz2lZWZf3zBoCrOC2KVg+6cdwaPI7g44h5eVpnzT6TmC
nXsvAuimhL4HCFUWT2E2W12bHe7zlOzoFngAhIwX9FJimEQGqdfjQsn4uGcTs9In
38AAlcF+AJ/7z5r6nSaHesVvu4iE+GrbB6Fo0nyDKLsSwC33BlxtpP44OY740gFE
2xNaegTmTjZdZmqX8xvJG7CARmVCXjNRP4UxT+aOZehkMpSDTd7uUJ6U8wmvnqyj
vT0EZA76fpC7UUVIPB3IihbYsSmHrMCwcVQF70Y+DDMeEGxzvSmu53sooIC97Ee0
MSBNHeDxrUp8r1rMbMqeQNEh6pClGdoDrGoy45Vg8ytc2O2sE8A8+5LJKiitriGl
xpzAT83IXW1XiYaKr1kO3SWDkTD2j75L6i3AQ/1THvc7ARvb6SkvvQccwABCmm75
VHl3ZFGqP489X+DqibCpRuhQv77w1om9TnZQIjyChEZTgHymtz4MN0JNr752vZHy
qjlImoVlmDkhF9H8AqA9weKEmsRtXF9ep3hMwhSdHzXdK8MghaFuTlc8l61qU6mP
NQm4fsTIYo5RCBgVS/oTMgtK6O3Y9atOaGz2A0xtSD5u6GvBhNMEsnPxBBshsbCI
NYplwrQ4KSq4YKG6+30IX9NrWv7uT6MtNDHWct7UGazeFtOPOJnlJhqHRh8V+TGe
jVh47jAVKj4CoJkTvsBzXdaFdlR+A7u0FGiFhmtJlzhpb+e+yLvz8qeiT90Ogcr8
vDMOjRDHtATs2RGkcpMfxrYDYNlynr5IT4aMs8VGvvUmb7XI8u5U30Xv9I2aaUTp
o/2MiyhS6gAF6/PSffRGpsMDDq2CFtoaAbrAKWPb5oXaMa15GAOJjCug2VdK0TXy
ADUiY/1wr3cyZEyilS3L4AuV0yibgemb6M3eu88iNql/CcUzn2pPJJGhCk17cqWV
8+bZmFSY3EOQUJ1ku2DNheAZCOva2xfEVeS83m0KXG82XaW+v3Hufk4nSZQXty2D
+ON2UlrTygF4pCAA8XZMwNKsjAYFQhqx8B+7KDXLVM/mwmt8KeR+RgQM3QTIM0XM
k7dnKSTHqLoZupUr1Ll5XYiL7TQ4yADqEABM5fuTr3RfteyhH3AYyPhogoq11AXB
aOIIPdDKZKZj7GMNbAOL+AAdYTHTSfLeZsDXjJ2WWI2gc03NRka+YeZbM0kpR4l7
kM0dlbA1vTxIC5DZg4z/RgpjbQEjrpsVnC0PoehOb2jB99yTIjNBY4Z1XnQNrZfh
nGj+KZR6S7wLfl0/5GD62hhlkjLBkIV3ccpJaDzA726r/WNPWxxgv9g1Ka5whng9
cb4MEc7GU8b+yuetHJMnKSk7f/7YNHb6T3GtHRZnkWsHih/lP5qBc4A50G7xv3q1
+FPMvK+QZMwxfsJ/RKtjapib2H1TjyMTOlYe0fNu2z+wNr2gup66rRm7ajc9aq5q
CxPYd7S+sf85K43uNkZAdydNhgGgTMNmHkI4Hhz8O0wRjfiKKc05QeQT4jP1Sy6Y
KuBN50Dv7BmFcCW2zD2AUJG9v1FRAI529agAy2Qti+syR1wIJwCiQiiArKjTgI91
1LxAZGzjeNQnWZ84zSYF9TqH7eP11Lcv+hxh/QtDhj8maDqQtiHLqCxroI1+GC1e
PYeGkQPIWBWjOsYRFAqy6Ntsk4Gthj2N0OeirGjMGxTBlp9hWNSXcD8WQ6jMriZW
whka6Af7Va2+y1jeLoZUcTNjf4EqJBsNOlGKgIRPRz6mwnVFJHPCmLkYbvfIqJyp
3IUHvrRkvyY8pjJ7aGhN8BBQQwbiLq8PXgg7TfT41uMLdjD4LywJ3AiqQmcYxcze
fnf4+7BjkxMN5OCguFMTRJBo3mZOQ179YSFdefg2th/FciBjzvCllwW4PnnRi1Qo
M0kb/molshFbW0yjmi/MenJDeStN15BhKOAR0p0cmOajYdV6j8DVfrjuBCaTDWcz
QFUK1b4X8+4Vy5GyzPUntJZ3ohrdskxB6cYppQy92wsfBqHjMTwHTNeKaHM4iLFT
Aq0M/kO/qBsd62K8PQzWoWN7qWbHCfZHUQ/tG8CQJEdIpScgRLl1x7W1gMMKkzUV
8C3tI4sNMGB98OGkPn/Y44lsKD6mgVbu+0L+E5zEn4keks0WR9LNok0ZnocWdgvl
xi0+jlY7OxSQxZElJFYWbwmWvLh8XeP4qc8RUra1VxHC9YWgPQCbk2zTHdvvJiPK
PadAAzy+CqNKrtkoDYMJVmBYDStCofg5hBTYJaRL6JtcMDB2qz2B6CWnskuDOWIb
y0cV3/TuOOKW7ApFhmIYPhiB7Yt/IKhFTv74gVmqWiawZ3oRdjRxZ+LnmGrNC+AC
hOyTJLvoV9yTLnEiV7iJA7cLRD3fDEmuOpLgdXxvMJOaRtACKwSQp7Wob+wWxVo+
fsWuDs+XgUUSAkCnwfptLnFGdkfPlmGz93T6manWCxzaq9r5+ehUsuwyXCekAZIA
CkHBgAYE10ebamI/PUsVwAeaAWxi0/ORoy3bYcxp765NrwWZm9VEcKdoJk+BJlUt
phCcUJykGvXOM/ORM3tvK7RrqxRmcRA7P1uVqQQFL2mX0OsCGwR4cIndcRWgwDes
W8hwcetJLtwj0eIL14krNLfuKUOxY1Y7ffmPYcPm8uke3p2+OaYOKTnQsqAa0Gmq
ykE8RAIhFKG3BEz9zrh4c44uRWhi1k0sHcDeLKxXdT1hAWfvAl0nKVM0Lzpa4wit
w3a/tExjIefMI+pzvS3Rq3NZa52dO48OCqWQv+4tuikcDK5cF0J8C8VHCqMXLdlj
CDMSsopWPHeE2Id/OOhLdxNlVbSPumi+V4tPy9D6say5ZKX03pHaqqFYlYf9aGoD
HNILLQ0w01e9qHHP2mEBbVDtyNuGttpEqZa6wCAUMI193Wleq15CjBW4Ty+49Oyj
qXSPMpFz5mGGydFOZskbG/GQxyTVh83MYEvT6b9js9Flh0MWbxkDT3xUSk1u0IqV
gat3FlJbBeya7e3ksDUSsRv2e0rnsOKHdAVWO1/dHJgokFh1gZz2HBc8bE1r5341
WZoTRghi1ldu1v/dJZdbf4v+p2l6fWQVUDbLblg5XEfO8TyJx6+v092YaNJ690QR
nYYFyuQB/Ax55b3VA0S6OFehoi4ZXXxuz4DRO7Zel23ZvwB+8O85K4VCAgytpVxi
CXpAM0wyTPHCz9Uhv2BZuvbRY17CpEYSHKppbx7GuL+/kTJLemSvPSQJ18OjcT+n
DohlOQWmvDcXCPLvpRpkzo6GA7/oFaYcqahGfQkpHAyE+IWUjm/pbThzETBEAXnY
5jMA57xuXgfkEagWx3KJrT74VgSwXivjwX3MmuIAT0W20jY6j/WsiypsBYG5aIxu
PHPB0Id2Ru4obIXEu7TdnMyS0tIo3/pv0NUQaCK7XyinlwF8711okVS3eQIgXqPE
eCU62Zulk9YFF+eCboIjY0bPCYNoKfnDpG408aP+AVMC/ayvGzJf05HxojJwcqVc
TofZBZwPMp4MBEXxNuP1B4DDXAkeUOWUQ1eADAFxh7v4HewhIbxlqZw0Xgcxx00f
8FuHspHVyutrMdW4/ZUsj15X+SV/vruCs7j8LNANL49Me8qQZ8o7B/sQsYE2LvKD
sGDN7LaIibznjnRozLl2xCDxNk6i8H3Uy+KDHd8RB7ButwDfRZ0cDvyG/W59n5cW
uf0NGTPsHZy87hba1n5w8E/Kl7ztI8prwheuYbxHKHvxtF0TuQl68X96DiBjGu/5
t5uFi2vjZiq4nxzLvDmeRpxFX0yD+QLMXtr1ElAYQhFqt2Ei0YnSjnHg+AKJn9Nx
/IjM3V3nucGWvYRtaGzwogOiwlCpMlLLTThB4ihyKLDocYhVaspnnbxODKCnoJyn
tg4rmOOMH2rMN3407MsMpPMgE80363KyPH+lCdfAqY9fNpfBcAvfCoVW8hpL79hs
qGn2gkRlwLFPDvJjFCemZk41cUknsDVvNfGdiKhbWFjhsf/5M0qPi0g3TbHYE0+z
3cCArx0aBtfIsBV8l+8bgY4kBkjEEme+9IWxAjLmQrGsFKRkRAk0ECsoRowBjNOd
jU2WF4v1P0IxISNhq3jUZPo9BhcfYFM3ZFFyEA/f1gB5VFkKcHZEvM1p/HpQNygN
VrXqfo0iNtgPR8npdVxHoTA9SIJeSWpmMCIu60cPVPSeX02wB2KLM+fJnSsuLmWP
KHPKHqltug03rX4ZCwYtriBEmwV75ge5jnGvsRgi+YmvSfBcWpGxlPxEyyFMT71I
2ZDgPQdSv6rCA8qi9dhvvLh3svWhNppnKwF+PTng0wcvIWsL9+r3E9aH44Y5H9yc
qBpW/4PKV6tXvlvHcjX22f8G5Bqej9P5TZwn5ZdzjAt7M20q9oQiReuqiETAXjiC
cbNTMNA4lB1r4GQdj+RgcBSMpkGo7TBELx7ZnIyFwEJVGHaXS+yZC9pCEEb+xPX2
FkD7o4vg45iynavf2pRCMc+48Y/ok9BxcoEVeHDA2lQoDnEyYq0EIA3zEHD6O8iO
LTk6JrnKLPKO0xQJRGu9sha5vxkyIT4KU7cNnKknFAqq9pajbYAjnYyS7/EbN8ut
MUh8O2y6uhv9TrgZFuUR4NUW7n3/LnPkFzoh1jp10pUhi0lVaDhAWqz6ycXcdm6e
EMSYxlBJywyrOrZCk3/sZZuCAKppZOib1PFaf/gMiDi3e7fnl0PJxaCDZZ7OdkkK
pPfKbz7Vjp7lLJdEbY2EqqtJp85hyHZPxyKsDBC9wHbkw0yLj+EYjy2iVF8rD5pJ
dn4Rc1FGqD124CSluSeHBy2bcYVa0d8Ib+2p3TDrKYsWkvYQzRmuQgI53RFzNGJ8
g0AEL4euc/mHK5JO/0UJYDMMmaqERxnhbZhuzHsN5c/BoQD4eTxmvWm233or4xks
saSXU++x0pMJBPsefJ2MaSLAI7U43NXnSrYSaDq9lPCRtRxis+/Hs9T25uiuDBmj
TVorUgv1oHsvqhL3/YmCEPIvsh1Q7mvJZnRp/Bx6Xq5F+G23pMrMj0lu2fLz7Iov
9FZukiy3OVeg+YyPBu3M91qoICNZ/+b/qY3J4zv19Ru2498FwsUB9FQ9bL0oXeP0
xLffw81vfUVVgdLhAvkNR0z4/OuGz9jMrw7eEcA573DWt85Of5POfcgrJfj0gg0z
SBXXQEBE9rNmL6WTYccaPD+XmtOlDnepYjNR4tXZ7jd1kvRX8Y71r91ZCO6w/8sy
WKzkkJd8pIEW3Ldc5dvFqeMMOtbDlJcp3jZ+TsA2bPLmhCiGcEhUjiWECp633SHe
4YT8D5DZ7v3xbzb4V4NG4q91SLcxVDB3Q2iPLFSRYZv6rNauv94WrzLfsvlpa6hT
CXkF7/qS4eBbaUVNr6l4GGh3iq06KzKnAs754ELH5OKoQ/kUVPdNp0Wu4ym9mAIB
x2TEzrwY/hZDBSr7Gm5Wm/JpmKQCMvD+PQxJQGWMVotkqYRJ6+cie5RNUGPPn+UP
E4bLjbpk4yMYBmyNkpzf4Bpq72LONkH1PJgA9IXhlKkwaaPU1EnVZBx3SebyyzPm
3Yq516X8zXBVstL09U4HWI3vG1Cx6+l7pxHepakG9VK/eEZTnaoO2iY4n0PhV1pv
SijkOrjuOAHlnY+p8o8zYxcS430ODTz6tCspHKElJYBPxaPKBfKp/PvGPryeYCiU
6qJTNFVmCP7/k66xdJh251m5JaYAxVcZunzkw1H8ZtttCitp8a+L2/jeuxJDURDF
FtsmRPMCPpPnBmWn+svQCANRc/eaVYk2JnA1h+tQ/w5ZrjjL2FFvP4C5lVQokpt9
arq0/1aGJZwxE6bEX8MxsBszcAj+d9nuy+7LjPvKBWMXK5oA6rdwdR4sF4au6etx
qUZrutrxHwiTEppr5miCsN4mV9VAdvGDQK8Gwf/z8qw8aKt41q869eDP3UkMPg4F
UhuerxenMfA89sn44byyLUQBcdR/BA23kY74Z6/LEhVyK9k5211XHYtHRxPWXxuS
lcTVgo4Is76n6jwsubSe+Ojacai7aQV3MZBGzf9P+it9rWRIB6y8AdmHfoHcvXbA
RaVh16rU4yqgs+7mj9mNYZbyYmESfiZ11wzrM++i6I97zkShw8gx7XALat5s6T7n
ChiAqTMyzPPOWBEqNMavSlY+IaGwQZoJFeIJrlXchZxOpkrA4BjvtML247RjBmG2
FJoEyTE3BM2JXoHdbFE+umSJTPIZJblw9j6x3zMYI9a9Yqe8UrFbbesz+aA9G/Gc
614uNi/BNpo7PzbSmcSijLIufjlWUT1L1LYAp6935nsq/gICEChP+XibXKOKUsnA
0t9r4kRYmv/7P8e7dbKNMRjpMDE0ib+pGjUmwBnIWFdn93sv6xWZt3y9YaC0cyW2
qJc/USWNC7rBnbmDNugC+hb589Hm6RJGm5a9ITYcCR5nLVNLJhVdnsH8PFGnocSl
+e+gnRptel+FY4ebIaOGsOa5WEojo1mPS/5t366fzj36AoGiS/OEZBAVW7Re4E9d
YjM5PfJCPHmv5sVFJIXZ2VPaoA4LpRksHgF0hQox8rTdT/7wEXXXMJbicnaVP2c+
Cfn26c9+K/YTHP9dgKADYPAYwHVYW6tqR6Zj3dQt660/D3g4YHThx3vSZXQQYI15
oDj5ykxcQYJT/OLpCMFYacGIRqN0P4t316Nz9lggckk8uA5FFmrGGXhqOXL2LEkZ
/s40ddZBPdajbZkKKLXzSYgVAH8G6XsYeYTnunaEymfvx1QVTF3j2Jy7N+oY2f04
`protect end_protected