`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 38000 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eislOGByxcl/gRn8UziAa+H
mjgbsd36EQO5Ail/O6Xu+bnFAm37taWcCGUvJOSBO6pjaV3b5vhpcAiUmowBsbMq
XdE7LJJ4p6OSXmZ0dBXmSRufot/g8baJ2Vwpd3EucS5Xrpklt9ZK/IY/dRt7g+Su
OInnRM6tpKcq1/Rm7Os+Zw9sn4DrOnChksowVFV2vk+VLxvrg69o8HNRU2/g8xUA
oYEbQ4CtTpREoQTagYiA1HpCz+XpdRsM4fVQVvzfGjJj1TjkceX+m9oZ3k8PkW21
rbQOkCxjDkzGc1KZh3h+FZyA0g6v0NUxVPjMC/r3Ac00imxGzpQ+CFAIfBaKne9J
8kVBifJ5t42lzxVeKBSNdzR0XqP60Y1FOci9LOiJG8zEkxcWNkimdQxfSJrfUK5r
DFzOGxTF4n0fI/r9SbGOU7IAhzQxsZQxTktbG+qwtGWg49eb+O/WXn/pPEi0ADll
vTSMexm6zoE9tSeVRylqitwnHJKBrD1OvsJ56kHZsCq1/gHXqkQ7ed8n7mTmIrdv
VeMTwJKFgfogS78xk6ZTCS2T0SLLpnliX8xZLoSS+AXtmsg4RIh0HG9v3JFiOZus
U9akhQzAy9VC/namALov18rkysD4oM4W6UPPSaISEKfP4qoDMrlxx1bl2tqjsj4e
ErqcfVhZmWde+Op/KKFpVw1JhkCx8HeisCTbcq2hCXjJoAXEXVvQWcOqubDT41Gb
SGUIUYdCDRLAwyailPvXraF80FGxWjUc31rRio2wT1nJ622Iur3QiUhBouxJX8co
LsxGfg9JXyRZgl7csnlvvrzSekd/6uJzzqCcXchz4BChbHV+cnaSEjjLy+8+XW3T
HQl0T6mBTckEEdxjc7OFTBYI5OjZ3WIeHrD1dN52wb5mofMzg0lvsYF5KGSfGCzt
eWN+CHQTj0CzDBSgUWmJ357X+zhqS9SmKEM03yIn+d1a+4JUHmZmm5t4exVx6/r+
NNgrT89GMLXVChi7lwns19cPMnEHD6zZMcADj5viPe4maQ53yM0OyQD0ujsPL4xn
bbRlY9KH5w1Dr/PlYXklSTnZ6bMGK8iw1//e6WQtjcMKD3PVWZqmAIZI2hztP7JG
vklPOxO0ROO0uJjdDWhiNHp6n8oslpUQo/70j7gaRBU9ClxgK8Q1E5rdLHPYinyP
na7UFyXjnKq4A4ywQMGqG0y1nVxszv+vLfs03iQWh9AG4XRSYdwdPId4sJ2/teM8
L9m2W1mtLCdK8epGrztQgAg00o3MGSB5kcgsyG3gEexx/ZwfxqUXsjHIjrTeC4qa
NowzMcqwKcRMzsH18ho/cSK6qM5r7DjQQULnQPon3Qq3fh7tomDU7DXxsSGa1P3H
PV7SnzifmssiHzOSyxpCSI2NpRAY3/Voh+kpvYAHTyDmm/0bZ2rcojmm7YCysy5h
xo4F1G5tBCtnMHouSQhdxe4sgKjRqJBRK9KMMBn3sfp0XGqZZD/VGtM09hq9+eaw
ifEtDfp6mBd4wqohzLRNMw+IO9zX3rAD+RN3de91H8erFo6WaDY7b7XNTnOV6ctA
T/V5QyYwwVfyG6Vb27V4Dk6hcWpoaf99XUzE7IKprL72nNxEANFHo0DQI8mX24bG
Pep6/LczBW0c+FepG/h1l5F5p2QxVuFmhD/oWVihbh2tKLPLwh6EyEBveq7q5N0a
RvGP2P1j5GSx3G8TpYRFP4Kfk5Q3EWMXV/qql1cHbyYOIGGshEd2+fBHdvB/hwK9
UdgbeJa+L2GnZt5piZ4MDUq+7w4lB5HdKzttXmuPpkGj+v/WmNrIeF58fBJG1rIS
1erxDU7pCdbLZYqvDb/D7+Bm6n1A5kj+Igj+ti5Qa0RCKQ5SjMw6xzM8uIOrqqfE
YyCzZKU2B2mtyxwZAhsEgaahr+aLZo/0BYpi046bVRbffblJyo+gQ95c6Lt7vKOc
t1ushunklTfiab5a/wvSHzpe3J5c7lrfNsDZ0twhiTLqUS+aNrKrISQtr9th3+mu
mku0KaTlzWcpall7TUquVyyjI72G4ZHPgLKq/PjbmoYQkK9mw/1sZzwXI9AsBdur
wJn2ziI36tkIAC5uALPuiuixlHzc9BOVn7jRxDAexmpDwW2eDE8zjfFXHKBTnB/I
Fkm9ft90i5KscR0BP1qPuZMGxjvJEThryBy3zJqRNQNokmGs5E4kOgX4rqkx+dqj
5iDgo946Qjjr6qowRld90D29C/rZTpsKDTfCWWofBaDMwt2HJKc9xk7PSm5EY2eN
6/Lb114USHHGQQh6zqbA1JC//sV9BjbE06qS9Yth5djRTLKrw1UmSAwHaXOMioM4
O948YI3+ByUEn539vzCdzrjgT79KTvXMM1gpuD39dv82hnMR2zKx6eWbZqMElBmH
0BAAHPKLLQswLsCdQhPzd8c0PByA/Js7nMcJ5nAfKEipPWZWKumjII6JaxC04xRP
1h3vAxP9OR+ckDuX5wvqlt6tfUMhduOZ9H7Z6X+d3EufLfGPe8JPNl8LQcU7jsip
Xir2X+PviBJR0M3KMoqrc3su1JasVUmixjKovOsx+o5kOU8HMUNGIzvANomqkgYc
2FoyjYEcGWwYf5CTUWwojEXa16gh7r7vqcNACx/csIHAk5kKP+07+XfqqwdKmlHX
SGZZajQf+Ueh8coy/dSHZpJ/8WsRYgUo66o9rm01C2RNlQg1QqHcI2enmGR0CC+V
5prHf/9dPPPl4OT56cnUhCGqczFKzKen0GXpnL8WHNjThEykxZShwdsXBhu9bDAA
KplkAtz6ctWKcej0hCSQmY0jgzs7zelqjBJhoIdmq2goACQlExztQpKS3B36nj7t
XNDdBjBxlNixxcrcuASIGfBt32yF2bJnAVvRzBvzJsZbB5F03ITgkMnabUG8YiPj
GmFU37+dRErSas1tc6ee7FdH9Kh88TCphj2LxUHj3TMNWRswbTk+hDKQSOg+QW59
YaekyiXhtp24GR3J14JtIdn1N6dfBTXoQx5SO9lcE5Wc+DkMMrNr0FtYZGufj5hg
FSGES8JU0LtGODYNn+HVffZkttikkDEHnUzlfTXW2zyYbyip926SgsbonUoLl2dR
A11WXSufm6Dt3kF6ig41eE/jYsaVvVIIJ3DvKggirDOjsjx2FfPv7eYv2zpwAtvf
8XvPhyCaPkZlR4KthiNRPmutbIVDui2oBPbaE6nECvi99934ABNPRMKf6zCNBjN1
plyG+lAuZBLp1hqWa+kNPNTftHDdMo3K81gThoJ6r2WDMH7NOb4+spLb2EFeSW42
CCCbdI6JDaKaCqSi0WC0A+yGGTyQIrj3txNdFG4ZV5Y/qvnz4yMlunIHUpZ1EiPr
s4bY6X8rD1Ttqhbwy7bUSbrNdE89AYvtAPhjjB0FrL8q8tTUJfSBGES4dLVKxXz0
d7Ro8Muek5Gn6rJdJankOAvltIGPDQGHISVtVFZv656Q3aT9KEozfPLSmVTU3VW4
zaC5RvURoaCfMrllkdxmJE/Oqo45kf/tbsqY0dg7KVdlAu2VAz2xe6Gp4R7RrQSR
ywSC8MgT+u+m4Ve9qznD1TZMWksOxGNqhCs4lQ1k/0WeGB1ZfmyfFJdIFzx3EaZF
epCMmNBkXj8gIH6h6rERws4XDEkaqsftpToS98hU7bB/JgOCjG2diZviA4uMvdGw
55HcqT+qCW1hnOkwbcetrCcjL9yj9AmZ2Wr1TYIfkTxB6ck3EVlQGaeojLcOeqT+
EerS89v4oc5T8Xlkij/n/yupv5BL17oMavGbTQZdhMssDsOHpp/grOPcjUHZN7cj
K/KCC7SWXZPDD5o656JdoRy42LRESeTXFBNWPyoe8ONKnE0opSDYy9zr25udK7ME
LwM6cXDFgaT0QaCPueB4NqwnOy+hnpc8EOW+55Mkb/VYvKjBTs+PQg6Q6tet2APx
HVzuh4hR6SEI+R5ECYachNuA1H53L7ixhKGbDZUA28zqQ60yqRzd1priIr7HbO/S
W4Qhc61q0CLw03u8h81suGBTrpUdAe2DQw0TKA4j7r/QaaohO0aYRmPoQqVqUasq
IVFlNYFQ16wiCFkvJHLML1xNyBNn3geHfJHNWGj2fvkS47LZUwAjrKn2CVfT9Gmm
cYHCG1NfGAzrjjKs7DUDt29sUCLFIFcd/VyW4PPa5b56gI4kCp6jpgGIKrSz5lYx
pv5kdw+XaoO6ZnLxz94eQslNaSuHVr8toXSJYHok91XplIy+qV1Wr1Jx0uYoVRye
P8bU9AVP9U0tRQHJGW15caj3FSa8hjOnqBRqnp6xCnKopMW9Tc22f7L5vh9TPbkV
VPjLI7XSLRV3tr68+jP1SNVkdFbZ+rkBQl9rznpABVl+lt8ITp8zsUvwqZJrQtgs
GphGhmNsHCwVPCrbmf27RnrQbGg7jtkdNip3L9iLHMAacA1zPKXDnpscPOAa0pGR
uPRYMHR3WVMb5tJsGiojziDCk7UgFsQHrVOvuIfhbNTjBh6I4FgBNQHLFVxnRUQZ
P7z7bH/Bi9Ut8Iomz2TOk4+EyTO1EKZmsvchs8tt/UeYdqJ7dtqX27fNrJs+G/kJ
ysEOVSZcVQ8Dlbmoj7qLMhzqL50qGG9sogenPKJjE7oziWOmjJqmp7KmSKf0v74M
YD2kb/DYkLUYr9VVLKXwBrFP75DIj6FBmXFJL0dMKvlNynpl+10n0yYUnznPZwzN
k+7vZZssvEfpZGXO4Ne31qcrXRCOztw/rkRnLssizRpmRtPFmyFhxzOLIjPoWKKf
oHEF0WltxVEAeSbLuzCPZHQaYrateZ27/nJ8Q7HPj8XjGm+nHT5SQKzMJOPsGt6a
yVCyyH1tzVkspjXDkB+R9Ia2NZyzbt9eZ4AGlTsWEUMzB6Fso8QDQVlRzly+8AT4
F+/QyIq7lpGLIK39TykvTbmr788lRQ2is1QZIeBU20izeq5j2HVUsFQGIFv5J+4E
ERtXwRRzbFn1rjIZLC4pKitPOyKH0YTgD2C30SEpYCetJTlkLgvGGw8QYmdWd/fA
Mi/4IeXJ9HVJGiCWbVDMz3K4uWzUbPTCrS7Az6PYVdDFM/mzrxpccbs1yKWS5Ct0
/4MqLo3kQjMIEZLR9NUtraBZcyMAnbRMTA7uBkUVsGlR85NeznA7CJN4TQOdk1CH
nl4uJ6G77sMfzs3zYp875KfVvDIK0SJTIEDrawuAG5n9/HYRUQnZ3xyigP9Zy8x/
5gaiZpK7CSWkRy1gsC5NlvtUQREIXhuXoPgMqwrLD2sz2i6CpE9WwACB3bi2TuwN
YRHPv5NGe4RT5cMmNXNqPbsVklgi8ua/pJi9PAdTcLKJcq3PtSie95F5GE/1/288
GtQShLao2/lHNvDrWhrmvL1qycuA2sCusJf7Tm42JrXd6OAJxA8E10nnysRVEvlC
uJZUyljtcnjjrFoNzegIaaV98x17OeZlnqXpF2zeNqCqs4gE/7mPonBTjenkInS4
TpGXMUaW0Rd00SUClNLt9fIIwWWysYGKZjrR4Kvz/zX+yaMcKVW2o1rKY+vLbxUy
QBfvMJcRMD1cd1ArXHp0EyqQ7YyPF6vcQ741a3ro95m65y63ZSpm/Vo9unkqK3H2
G6zYF0S4fKDACwV50xzVquJ5ENSBiM99zxup+U6wRnLa0KxhzbLzAWw+QXbrGNJ8
NFveBKI8e9d3LPRuT9Vu5BjAHQCURxOv/L6SK68TrnyiafFZurcaJlFIvEnFO6ti
xqMcL55JLVncgmYyQP9LAmcGNRdvxjajxIywewt91sWHeNlJII1b3WvcUUK+EH3h
kAgp54wIKCL0hOBaOBdpWculOJbOjomeameDgE5bM4vkWmXqnLqCXjNXlrO5gT11
Sxhv/csm2F6Jn+Ntknvw++x+DGqYBbkK+FAT44k4mrNBus8oKwxzjJ3CeZ9exhg4
MJldPBQXyyciRHz2Hie4o4qFqkpD16Twq8vIwbI3iXdZveaIwlf8GQfLLcvj4R47
Kwgo2OX7quGwmHnkLzVEI3eQXfxjLzL03u7Sonujj9m6ZfN1vJluwsw9NxSEVstv
SB0SvXaLOm4ycyL7I/nBOUUqytWkUoyZUx6c4MN7YDPdj7NafX6JFEgXQXPtMM2L
+OwhekD45ld/Fx915CK0h2foA3YH3LFKfuh1aKe8UXECvOHmK5KXFX7SVszF/DDu
90Fr1okpUmWETfuAHSb04HLDwQST8AEooAoP51JAtSRUKaefPQmxp5prOp/IQaQC
6UL7mtnCafH8VR9TTtvY+7vOQLSCC1ps19r/MClvoECSY6MYzo/otJ/HN9LdRSPB
JiLQ7cxNKvZRCWqqOGBDROyGxmInnwNFCE5RcVMAgW3QSDrlfMdFv2k8Zp6m92JG
3eGBe7A7XqQH8Jr/YTrwf466od2jjzAlcfowEVFQ45rOocZAaJ7XdhR8goYxGqhL
yBjy+4qAWq/OMzABHYvipGioMLaCoVpe1GZNnB5e2d1a1Sl2ReHpzlkrgle7bCqY
BTgnZxtns/jZN6kRAIPJtXNGHOqjZr6EUBuiokHRRHHC7Otty/p9+KFFN5CZhSz1
WwDRdb6Qpvk7EHyXhf4llZMTagNbd/hj12OWetg1fDpwcEBzQxsgOMbRCe6rgMmt
3xwtA0hJjiqtJjgC5c73kLQvxEl8sJ9y908UcDGC5CfdBcgPgBa6KLjp4FxqAxAK
9s6SiRpJ+myGg6IjzyVKbYIBnC7fbJ71l0gm9c1z4lNdosYsjeXVzUDsYT63pKCa
3Qo5AlRV6+QBYUmhUA2nbAyidaoRnbRgCDWvK3mKNstd+sNEiwCm95g6/nQKVSdE
w419iZG+GpinCJA6dWmXMvB8b7fwZMvrvvvGp8DC8nqjCGxn/5XudUilDq5GC/aC
TJftjCi0sHsirkqw6mxXqa3ylcHFUICPr4YAiV6fWjVrru1Xfcqx77bF2a6krFgJ
3Ml46kHqkFkNelqtZGv2tG6g4ZytY2z4n4NZXKOScwwyTjqptER/kJqgqDsme8E4
KExs13nRNozyWGMF7WUARYQRln4nfX00tpLJuZTqJKkvlC18J1DxhTsI5UoM8v9B
HNFnKJtVnHRyL/i3VjMd/Sr5to+/mDh73UkuKUxz/HKqaE+msBMV84zX9O/U9M4W
2SP+c7X9aNIZnO7XMu81m9tcEv6Wrxg5FnjQTQxuUXipWBMeA6IZEC7lyWW/QXzy
zoPUEluMGXhlPVT6omk53YPhzDOsxt89X8d/Z/I4LYliVFm6KGn9aK2ZjHMWcgHh
O4QEn4UFWais0V5pW5fy8YbKsrWSK+vhCizTKsIs/VO0pOI7oEsVB51/1BGQpwkJ
GZfuMfWSiXHqsSM39lYXUNDuBK2KkfKewAsXDzRGig5Y1rB4XuUDjlCMzE6IJmFb
gzOpNBhtdzEusIJ0Qe4Sk1Xcr1gh1z0cRRMGMuaRUNIm71GiHGYBgwCS6pIsb40Y
uQL/xmmXIb8+U3026Wb4QNMT4qViw5hflPunykygx9wBW73HtKMF2ZTV5LHY8oWV
BRQiy5QoGzXvbkiwJYRqyWEuP9l6iX3yFKZUgqa8RxwCommDOFWLkv2ZhgLLSXuw
OgwDczCdjthnoAPkeMLjaR1ZfaZX0DFOXIvu6fzqZR9b7JPdH9AKrAUS3ix5kHXE
hZ06SeeU7wWYxaMgH9G6ZzW6R2PI53U6a53tG5Du3wUZKrMuzMDZlb5OSmiyTfX4
Zvk0ObBMdeJ5H5HN/Unowfm1rv5zNEGRLaXg2+a2UxXly0bUf2Y5YaaLz+dcUsex
8ZwsTJOy836DBvJJSQ60yPg3Pl+cnymMGt1glBBkvkq1lhyrKUBYKWXp3i+8M5zO
q2ZO0BsAdPc34ZrLx3GwA5FrqELaqCO/okaPU3rHZuztPJ40SKn5ho6bPOuIIj2J
lPa2UT+dVuTs8yYhJ7GD/bP3rMYPEsMs+sQ+MInatVNgv3Dwx40khOll0mtzJDv+
wuZ5HwyuS/y/hqQOiEXftThBaiiMGj1A9WgW2fZ2g/GBxi6CNGCmRETXjfar5MRY
rSu7xZAiT3CLrSsNMKvSMrbcmtsKmubgVFmAU/yBUzyBIjbksvJdxaNcckaNjyud
ABdAn0jKwttAeQARJFC3c3vRAuUV30/HafVYMraZFmaBvPcrKvmgDXFD1x0dHvIy
rnVmRW7pmH5Ah11dzQZjBc4/AlKRY6moSWnC43YSmcy2+rF0OSxOJFrvmb5ksh8H
Uag8kgWKrxAakj+aLJzSiOzCPDMTpQDI+3V+nLpfhFPv3GytgtddQPjeviaJlyu9
8EchxCOIJs78IgvypDmxyx+Py1oteiyT5bpMGGBn7SCxMirZ+v9wKwdrPQ4SYVCg
x6kjSAnIbc1fElTDwPCXXktQGa33lVPKFU/0rYnynvOWubg6jLASeInb4mt2Xqsa
kY1B1nyay3aW6PCln6w0rdk2f/mW0QBLkctWBlvzkWReisOKUvFYO8IAgNOKQ19g
4mdnCRfJGk9DkxR/xiZ0nStvd3CtmbF+1HjhAOF1rXCIR8+S0pNnfzyOjV55CkQC
GpSf72HRcyQyH75hUsBHexHDwwpPcXQTFt31Nwy+tazdkOcExrLECwAW7x6tONox
qdsoMv1HRO9GBe5+l5KXLgH4XH0XDZx9+VBbgb/H4JICDlL+Of2nPjjwkgASbjmJ
8rg0LqWYdc2QL/9HBmL4hxghtHbuQQxIn3AMqK9Am8wkcNSR/yhP4sbwloQpwJuF
x2WnZYGhFDjIpVC8o0lhkV8CfNegnZ5lCdnDh5DxfWpHoi2N5QHlOcobwC5e9ZNK
EriDTWbeM881E22m6hoQp8qq5huxBmfZ/F49hlsiRbhOfhl7zY3+xOYwyPn+pClq
eEcEIADCZTgs0CLj56LrkkrXtiCVpcrwAriIl5hzsmbKkgouL/VxJNgdKJUef8ju
d1lhQNv8e1BD8VhhMjXD0BmIAOQa2R1PRUCvub5CaTEtLRXmbiQI3GvtBcFsHgNS
zNtFpBgwwEUBPS66YFQdfAJdmqDicVzN1IzBWZGJEYoq2gWtx9BozzO2IRtHy2Ek
GhLoaJAW4lV3qeYB69tpwWHuKUZQXuTwb9SBO4j4+p1IcmDBcxuoCm9dxpmzsi4+
bSYzTzwkdtwLPNVN7h8gs8GOGioBVhz+YmYvVPjRVRNzBWyO+9vOYNF4EK764XWL
jn4CGcXUuo5Bm6GPvIARKUYdm757XClTShtQY8qzj8O4B0zkRZbUdBMu/M8BzeBL
E72gG8+Zbjws80uomqnD1RJQ4wQzDHR+qduoRC9/s6YDmotDSDps/7fvX2D2pyqf
CwsIEtRDsBz/9r7uoqpCyjT1BlmxbMGDqynS/qvKMGmx06y7KCWzlELHU61vZazO
MN2ZKwAJAhVnCqio3f1Q6BVnD9R+7lzjXN3+jURl1kSivZcs3y6OdXpxoHyq20ho
oeJRDroLKhbUONnid113dQD83+bOd2tyMl2WpTR+oOuwXmqojhnoEv90LCaW/OML
O0ChfuuyP4/A+Ji8l1xdoI47H1cD558IpyaX0yyqyqH5NOna88PrgujYRq8Bw5lW
edL4YSNUEMfpGmBtweisUd8ysYBT/vs7kViGx8cgM81fChZpnrYPBlsoYTs9Ost6
T1Su36cS8ja1cedlewuLm1ACZ0w2AtObUCy6abxImzknovGIcyTvnwawWYVXnUEG
9npxxLeVJNLLe4Ro8Gl9GmVjK6bGbpyGOE7l0yE5deEAjwM2EenksRHSXb2mZuQV
S9nkVOHomk/6NpaBzsjE9Xjgq7b3oByJY2zhxeCdLWXXn/b0Fro2OyaoydZ0enqs
G210mmJMFVVna4RfqVmEN6i0FIgahd7pszuSp7++wmjtQzKueSbnyeOjXxXn5SC9
AjFMwCgNfwSnnMlwXfWn7fg+uVzGW5Ki/4VBBitBAAkqLmRObYgb52+JcYY+0Ulo
hNCeNcNUBZNQ39jdQRDFcmMfVzUVB0MW8j0z94CvQiSMiil6OIK9acIDrineh2y0
qwd35XO/BnWLJvZDJ1FJeWTPZN5MK5xHHgQSGZs4Rv8JLyOeYpJHQhkxWxTlC41Z
xi2TUVLc1HO7jq27bqYK69gXFcZv1c71E7Et1lr0hY6L7ItuZI2K69vfWEhTVBkf
1l6W0slCXo6mYNDGvDQjQUW97iXmux9SgzrzFPPcmJfk7JaDNrWLV3gzyULshhMZ
DsGsaac1Z5LAp3go56fDXsyKxvIA4/gWo5PWm3qlqPfxvxqkYUut/7Mfi4+az8n/
uvrHTShBZv+aCT/KvSmvYGaOMVK22TpWep4sJeshoNNskAYemJjO1r1vvC4/Covd
TUXXM3apDFEXVpeMcRVYPzZss85i8sjlmFCQgjU2IYOE07ml1hB+mgLGGbuVu6ZV
rvhlNAqkMK5P//JQr0sDGnVrZ1fDyM+ZakhxZIWM4HV3tlx7sCjZmPY9nPLJBpi6
trsXieS4ipfc7WFDHaitKnrDzkarWufOsua8mgTHSgwzfRpA1jEey3+MojxXV2P1
r0M054xsnaKiIiWC5rM+X2QqamtuTgfclOsb2/HDoT/hwrCue1YN7xxwV+Botd7O
o17W18aL5SLRjSXHBQJo6bDZ0NdGBCfbxf/3k6+/YCTXMMJg8acC+PoS00EVt9ZI
z7jxIpWtMzfEJXEb9Jau2t2cR7lchk+De7E/pE+T9z0MK0aQRJSCYy9Kci1HWepM
+klZd6eZqf8MmYD/5C9VJWOS4mPbNPCAXSF6X0LccNBD8coV5if5ot3ulvEfkO8s
xdtiBnr6Oz7lmpYPGD/kQ1AJdJWqzhGuHIpsfvT6MVFqYj0LPHnlwA8M3QgAON92
hWgSlwIri6bhENVdLeme8jOTmlBvrb3VXgckDHfGqlhgritaLZkx5DOKEynyXlIn
T9pGmSq4Iwvy14REzOEBafhhcPvT5Q+hsA4A6eF9omDvecVfBh0/zj068HvBQw3F
eEJrAFjTdoRm9yN4V3qC9nMIevIcvis9rQQIbiMLm5p+tGgnKoJtQIuBcxZrxrYG
C/bPz7bgqNhtJdW5rsgg93RPO1AodR/4maw4zCizTfSgyISLhr+7SUveRrSNx2z9
iaQ3Y3Bevy9gHvujFsB755sGJrNQBaDc/XXFElM9azSCmh20DY/E8+/xVnxC8MKk
/xlTfEo9JS49deTN48rMLg1gYgruwbdoMSW9k5eFR9A/mZiuZPVBm4sjV7110pX2
uv3mRcmHuocQLK4OHbaOC1Mvk2IV5wodXb6K0jnaBmmv+Qdx1EqOw1ucougUtm+X
IcD3qRX4eAx35qmnEew0iFG/Dx6WedlxbQ8mzkNKORZ8Eusb0ueP1QDdX/TZCKow
xborvt3F59QcrzOzSdngopcJFkU2meNupxSpgarfOLLLyuRUi3rpZcZW6jdIyV96
S8AlcVfaPCLyC7kVfkUGFeUNJTTyldcFKoArOjyg6ykEmtlBPEeBEKWBL85jsact
7JUwGSa1pLyW+svIbITQdR+4Y9/0n7OeKR5IuOxtbqNe41vDbWKtuphN8N/HcVOS
09ZvKHY9LTeZgalmDoG/R9f27MVKOG2DE3UYnI3R2g+yKZaqqp+cyPhxLa+xtCvr
qB0WmvKv7NhPZeQ74VON5zcen89oBrx+A4wxkdC4K0/aUyOnjTSx6bX0+hd+X1g2
Eweq/2CeVyCVGWNC2cwmzgEiKKrM95+9rJN5KNZ4HbWPyC8/P6MvG+rxCHz7KDKQ
CnacTudUmfB2lRu/FtADrLfeipgDP4w1wyTedxJE8tzlVLZdM4oYyjnZZysylZL+
trh8gJxllsj1EMD9OeMZ23TXFPzOgl5ayPU/OldLZJ73B/OTHDbuqcn4zi3UIUBa
GZyW/bxMp0RIDtaGTzQb/7I4hKjaobjZhOCI+N0cVD1zgeBoNFa2L1hCvyWSpknu
K3oHxlD4NgrfEtzdvPtNed97TLhGE4cjBCPJBMJ2y8iNRMX60sYLIhsACstG3C1J
uwPVLSR2bz9bZG7N2BEOBkXZfdqKwLjCXoAV6n117FMiyW6/gPAenTGeE0E9uSwL
pR3MkYL/kbJwSUgRQrKL+vJW5ZF83sofx2+GvIqF06dlNu8sbdKXMr6JmnJNuffA
9TsLjFOdFOb9ObifKeE1fZFpiAh/3sz+resXQbgsz9uhjSR3Cjm8JxSu/YcRwfjn
N4F4Z3Uz/2yD78aNzDZBybzKy5oFJWLwvkaouhJ64TtywIqiMqSxkr0qoF4+NNAD
8r3j0veDTOa/pBd94KqlXfDc4+MfBJZ0xDYFbNSykux5gpLz6ZalppbfeL2dYWKQ
ufOYYD9al4Awde8NwLhq4izmQcOiCrBmg18RJ0dazVSvKtA3ZxXHWli2VkWcNA2I
VqRYloN0JOirp0FhKvy1IYzgnCA1liI/xMpN47nUQKmuMHsz9nzSErcJtpcP+Zih
t0DTri5O92NPMI7F5nd4RVuAEFC0+c5wbbvwph/SME81IL48s/Rffz4P/qi9psH3
RoM5+cyCzUn+RGbtMp0q8l98TbWjMhxo/81weYcSxIYwMTp+ULO7B6i42dYPxRp/
r5uzPIALTfekDj+mlEZnHipqEqEspdLXrSDLSuu43JIrw0qPrBpeYCKgklrwDYdH
vHHFrKhXNzfbAonSy/F0xzCtv8YwoQOAbmEJ/ArCkpJS1qjJ17ipmg9bfZgNkpFi
RUjZFusY0KwXZmavqQL5oLPksjQo+qBZHP5dIE8XI3iBTOQdXRFGrMR5cS2giD1r
Vo63HEbW+kybz/eFWqNBKsOMcwa4apytMuWQVIh1tjHGUQgnNIXRxedM/F7Ln27h
PUEpl8LIDwGeqzB22Z7BuBwwSIkiME8hSZvh+LzUljOPKX75L70Ewt8ULNE0TGTF
rDdHOeTsT2Hz7UX0C/i8V2v4//jG3MJ7SSPbUgTNe6lYuXx8cmIBN7ZZ1iFKUVJi
U1YRbSTiGJbugxBCaygQCJFoXcISOPMyujyx7aHfufX+tIOQwQ100VVrECHW1tZV
qTv50sP/DqpVkHaUgA5AUIKqDEnESDflZ7Q0u5jD8KVu4n+xs8toHpIpToHBXK/v
pnMnV6STwBaK6t6zVjdXbIk6h2mc33h0cmbRhFNRhrxvmBaLOVpH/JV9c6/pAeeW
7RQrSTd3ogb6w8/lL/HQUkW3/6uAME3Mj6HPjWTB4r2MJXgATRb+8WOXb0qWRO/Y
/wRuz+UqyacLCEVmHrNUyTDN8XqKbvc7vyd2E5H0IklW/03b2qNqox3a7+ZJOtdU
e0avphLU63W0L5hxIhgqER3JQzDNkR703gJFDByre89x7aUhcrGvW8XlZ+SUAhis
rq/PiaZDZp3R2Vk1ds3eJ2O1VcoBaLlPBHZhRyoaZzw97qdn6Wbme1MpFzY/9jwn
86pS/QOKU5rXh1G+/zFwZNytnbBnIsaICTE3YDGWMIQxMo7SYqGMFUfmVizMeNJM
SRnxLn+K7n3WMHFedjFem8zEcisKP8tgwmkr75sJ13CMXvbWsCkIpGOcyIaIhAOo
Zm+jq+K2RYdiW326ZOd3ynvxoSj7YJpYebBaO65cKjRkcKsTUqJ2LTtzS+xhvXFH
0cK/HyaHFaAz0PMfbmm0su5yhwJbwGH0+Czty/g81VieEGtMN10En7A6u9ZDFRNr
L/CQbIwH6oo9QGyfDgZvo5rEwEVexCTyMHbZvM0kOU4j4AdPSJurMg1hV2Wddg5C
Xo2nHQMEdQLZQpEztxspqaSfZW5IuTVlOU6Sf0IZyDJxV44UlgqWlItRExdOD79G
V9iInECiw72TW2wRJF67RwnlpRHYqtz0Y9oVauVQCYrV6ZlRF47AHLd9gfPvwGHK
mbe4kMxsPrEt0t0IX7qBc251CC8CEpzuNxk/HuNBPpzxq92FwbTr3dm1/J6h3kSo
AMwTAnV1rIGI5gWOAAjttqi+kWR6MJESMDbPKY0PD4Y+NTNt0FiVZXT+ZbfCVSAW
4j80sqZT3Y/fl97rUCs3Brzbdh6Q6M++atiwIEvAiCnFGa4CNy7HbhhE8ddD/ilI
sGrza1GjDA7dcFKit6u0sDkfwa6UrgJPWmuhMnAc5nBDgxXBE0/NHpmgC8U8xI8Z
fqTaTHSv9fC67Cn0Yi31oO47CXcKsqRckQgAHhJ3dh2ujZFbPT+p2nd2MquMEEKV
BtziwhhvUNdap2vH7qnwTjAYn8JDFHkziMwxhLvoKBnCWC8izflBKyJ+xKnJ3s40
DgxmCrwDjkgtN+/bxJ30k1fvQWBUm+iq+n9VIY/N3d9UdTFcHtlysKiWi+SLNY3D
3hb2IVjWGuOfDgGFoE89n5mburTi2DLoFbFE8bjpHRy8js7AiwkaxlOJhs0MRt3c
jSqiO5i4hjPmsLogDg7t8FaYXCL0hsmbF3+QiaUr/nYHqMJYQb8KQveKl/nJXOmV
C87TW6rdDlgSJNtt/zrBlGVb2WVy2hA6cwV38zSdOf/58UO1FRS4W/KOGYT5CQIy
RrYKWQAUQKP7yoUZNJoBOVs6Ws895eBkEwNEGRzSke/UYJ8rBgu9CBpAqj+4gPu7
I3E6pwofHj+SFDvUOcbHcjZ57Pt0Oxhcr9q9tOMlEDzbTOnvioFuc9BjlNGV9aAa
JzUB3w4BefAQC8UHIdr5X+NKLRdSC2xsRTZNm556wKzBgv4D7h8rh/yVdhwrVVxR
wOUdDrMLOOCHipgw7wy4dyLyFQaFS+3kir2M+NFowXI0Nthq8hmFOH1RvcUrgseX
sZpEUXdXJRKz4+FK3XsoTkKtSgKOz/l2uP6GtmrcsvbjSVz3ZCAPHoXATcoSxziA
9r1AwHWutiCxa6jnR83u1a3BcltcUrX/imxR9EKzmzlwHL7M+7hU+8dwx1wVWcIz
y6ppcvASZxYkOqRRPSsRMaWBly/iOtMtYBEodsjRxnSsc8B496ce1RTja/vgruyu
sTqtIQNctVxrnex4h8xxKB7daXcG2B7bhI8np4D9OCAnwg2lGhCsle3tX0Y9PxiW
aHX4UffAwNnMT16Gzm/yiKjwHlcerRvZIRn77gkHJ/6/6zBMBGhWu2PWWbmFrujH
roD2QfLW6zXgMrlojL3KbnUlgH+v5XhT3EtIE+4gXXXME/+/4rPRFaH0+tBLmiUM
fiLVmpdCx2iLOB6OvkcEk7Yhqrf4Q/dNIaqkzgQW9rid45Yq1uJs3G/LhCVYOJ7A
nrM2Q08x5/JrYwM4ZhZ79tZYcI411WwrtGOjKfvUF1wL8JFagkfQ1djeu5NnlTH8
NluIl2+0E2FN27eWjAuCiqLypckl+rJLtJdYpi3te7GT6wQnoIR33NHf8jWwKhUJ
nw6SfexBPORUu9luehDHTyKUD02Z+0x8es6b92d3Ku1BAV7+ChAnza4qf/dydm20
hla5x90NDGh9KN2UMcsEJ3rQe4Ioy12Jop/pqXFpND0LwRbx+nYU5dVbACsYbj9+
lfAipO5gyjLJb4GR7ciG/tgOaoBWp2+PBqSlHmOFFVlASXtVeVfAgITDpFBpVCG1
ybFOAvL0Pq2qAk+sPRyi8YIEp/3rSkMdeF4/aIUW11sl/5izV9QTQ7F4BTDGSNue
U3ZHMR/t4fVeBkke0EdB4jNzfgL0FOdHpQei79sSm94tV3JM6FyVm6Ix/rBA5Mm+
s3rQgmxdpcBYt1HPGiCcWbNoMfWCc0tU374nMCYWLfauUD+G3UaOp4JlsZQcnjEF
SO/XeORv7QlQ6kpM5O20NDXWpan7he7Md69Xp830+VttTRGb/7dfrcjaxH9Ab6ba
V2ZWPIlggTvP/U84JUxejtg0Gcx3udV2UFDO8ZaPurzvQFe56uPxpXFjtxUl1R9D
XaMbmm2s1oIRKLU/7YnX4AyiNG7W+8aoswptqPbGwHsM5J9CQdJCgMXdPRHyQBjd
CAb5yNpwLB2iXyes+f0oTAR/QwUsPkPyaUs3keuNbEcy7B4pp+2byd2uBIe87iBg
oTSBt5i/035SRhQ+igIH8FlNLKebejuWXvWKukNMoJ0YfjbPwx6xTYb9j9JQEjQ0
ywI7qB3GsQeP7hIkM9IeJnxXRQhEYb27NQV+TinrN7/4+310IEVr/k8rkcSmRKld
aiPGtpYz5dFW+3jzhBw3aqYAq2y/gh3ilJxvYjTVbK+VhcYeg40s635thiT9N71R
MQ320EmeNpQ7ihT4bPFiJuZHNE5gFcjIcr3jPuPy0dviSApDKNWXYoh5+W0P+aJu
yAuvdzkZtsanmPbwonGAf4pV8wkC52ycmELqX0/71eWM0e9qtm0X2OOxPOaZoro/
8FHHsWV2KELGz68xIe9NS41T6e6HfYjK44mzSugUEcYyLwwer+Oz+m7GLKvUozFU
JqnpOsOk8AS6IlOS376Uj5DnLtM5tVAotXdt6gziRZYYEER5edIJZHCtsotsB2K9
L8wvHpodhVVSDCrozY4yb7rXdgRcbkPcNF+fy1fARaqLlUIexER2EMkn0chP4X8U
lZiKv/55CiIkjZnE92qK5S8ncG/0ygc7gifgLlVYkACtiXQSyfHhssF9vZ3S+XKd
Y+tohPqhtz2AfZJ6j1VpmuWPFCboNPwYBEHCWLwqzckz+NpALxH3LsTbULWfiNuK
u6rei/2sy6tQKRGNmeje0Bl9kHueLcr6ZyXZLReKfx957F5gP/J7cTb6QHOAfdkN
7LjbRJWygXZu85NdGIGt+yTzCE7sjSt3aPqqw06HSjk6SY28wfX5ZF5R5TbaLobl
eJMBqsBdb4mSm/O4c3hbwlETpAH/Vx16vq/plF+F+uYq+vgfHT0iSdCs6mzjtsGx
LASegHmYFaTaPVvSeL2qHUCkYbLzk0MlL+WRsrLySJ0IgBttpTVpLYM2XxZCfIji
12wUI/UW9ub46OyIED/XFta+7x3sEP7n2up/rIbAwC2I+tWOKpJaCXn2z1aV+WWJ
TieLw4Ot/Bdc0jygbBqz+jO0YRx1SNrx//P+9YMN6iu7qoOq7UPfJFua2yF8vTVJ
1lQOEsYj7P5gvnWhvVtxqoBgoQjLBBIgBUsU9KzjlhyTAhPzD9TSkwoNifP9oM4Q
2nYCF4GfoMVYgyLqRvP1eLRWvSPh93O8IbsAU4qZGGgpAMPFptQJQcNfVVIJTW5h
Nm+f6u9fiCFwouWAWw0pSakSr/0QDlwDyFtruXc+KzHdVLmeTCXVStYC39WbVBqR
W2SOtDKPPXcdaPk/aDwiS3OG2Tfg0R+kY+Ifs/KMNTMlE4hzRyAhww1yuFBuGx+r
q1Z00uq6MeNIy9qIIb3/ZkzocWydYKzZ7rjpvEG3nviLcCAeTMNkve7FWoSU2BOy
ajgxt1Gd+d0JeySJRdp9eGImLZFnTtI7y2QO0wc9VRNnVHnh1cpGGjdiL95j3OXZ
RENTc8fDzb7c3Kcg4aXbjsBu9BxjHJJaOcRLQc/EbM7N2lrV3JtzxDhm+ZypQwcX
lMgYn3LUkzSXB0063v8llxkzn2veVH/Gtus9oGs3yOa2i3iyZPQwuxY/iVRJVBER
L0M+o5LPGv7Wn2QkSVLRYUJyZBj870qMGGF5w0Xm0/qlbKjnfX5FbE1x5KcnnoSg
EhR1hwWOwyHCRumXMwvMkEKfDFFqSK+7ON9ihrws6y/wNpNOsUUs2HD9XN1QKcz4
gyp/vgvsjuPUUTJlzO7tvmg5rLDbHNww0uCIWXhyWzO3KyKdBP0kG2mC1eHhu4Q9
LNVzx7Xl+adKvfa1KpqwEHwemCcAJVmSQdwT4AM0OIVPJkzK/IyZUhH+GvpE3ajG
KxjJ5pwquaaEz9NrdQ89rcd2UWQZnOkPOJYfSPWNeheHFlp7Ao3VcFLu+HSZ6tVm
fb2R+DhUSH1IR9PtR9qQ1G4Dunyr8JXHJ3Adkty6gqGRsHgGg9lr2C/n767ynpJX
Fr7z8zFMc8KynyiF6hGUiaLQ0i2roZlP7WOyvHLUJhzJNgjzvXLLc8oI4xxw9B+Q
2MqNv9SZuOxYvTU06or2SfCCUj4WKx90o8PJ6xEOrxbtPirU3C0+ho12jxNYV0F/
laxcAOIIfHJqcclZIXoN5iUlyye2LupblJyObSn/9qCPoFAjfL/efvMm0vwFyOV0
oajVGooPR1WWGZG+4DDEvU0UPho08Mnwxnm5ncb/pnO8Ci2HAyKIwWKfVJui+JuB
ZYpnYAoUnxgLLn5y6OYnVC4ynMed7hbC+B7xvb6q+yvVoTmrtmWvUZHOaVFIqxHA
MySGB+fF7GzenTJS3UePrGNUK+aSwzVbAy75rrlEngJMPoqn9xxWSsTcuyKEo4G4
+XykO6eAa53QsSZTJgtBKkUBiObtVjyb8Nnd6AheJmUI/NjXZmFjje4cdksIcUut
kR5ww64jmCql8dreQz5VzuDZTSvrgU9fCLtsAbPBfyStvvoNkU03FUJYhogSciuD
gFp/Vm9TiUrhyT5dWRaRxgyhwZdsollnCMu0MlfNLGqHZyBBGpu8LPONGvW6Q+3m
51/tybZ/zDVOsV6/b/thsPHRsWINXmZT+jLXkC3N1nxmPhU4j70wZtx6oHRCubwJ
Eua7dofHQNviYLMyZKBPoBeK2AmWQLLfqXavbYH5Yl9yosHVKviZaUywo5HeQo1i
DN0P5eq5dl/UVmw8ZMelbrSg9flRrQveRZ0wuB905mfBv7Z+KHChGAAYqvYi+ZZY
7FHVL3yDwqwpNZsO3TY9sBmyb4fmUP/I3MKgjxNwOEISM7CgmnpMVtX3fZtvwxsb
Tyeqqls0j6zVfiGePQMTOSnKAzsT42VN0HaNxx5fBmeWg3//NEDFWsqE3QC9FUoy
jODvwXuOGEhfhgdDBmNNAdfgSvy3FgvgcFgviFnke8M22SBI/O2rrJJEocADR5TB
amwpA0B4dHZvdd7b+V8oE7aXsRzdKcvSNLezLanJJUF0Yb1GUqTRisxD4HhphYbp
BjtEkhpVrAfu2SrzE3TKgyB7gYZYJZoYudr+o1hir+9Mz4EToW24swTF69V1cJhw
JwipHvv03/K8K3dwJumQOrf9mVsOQEYEBhEz6j33coSN6dEpJzK3P9X5QgdxubRT
E8mdIHxvwKQ8t1xLMesA7wBbM+aBxCzbB+suH0Ukjqt6UuNaHz1CiriUbn+r69FV
5/xl/2urKce7ifi8djElfXk5JL1UqdNQwl6zIGFRebWpxqGMpBpJScCtpDpbMszi
wCnQOV5czxfUGhpS7GFsXLVDC4suDSms9uJqgDaGUWiOHC0++PsMJYnMTF81UDib
Gqn+0TFGy/b+bhXhg6Qdne402xsY8k54mOR3j4amITZqRdpLfplMjz9bZELNoO4O
odtB5vXRpBKYjJjxVAvm1Zt4LRQiRxTrlz0yUfl5C8NFiMp3E0DVOE8IvKz1qgIh
NawHd7W1Jk7L2qU9XvNZQpykOT4VnxkpK4d4HHepukYztSWCFUqIwDES7dAb0bRE
1pXMo33Q/zswo1Ot+SO57aZ1aYzoMXs/VpYZluYFpD22zBYrAvQ95YWAFyCT8Aab
B2xjNokdiruc6Ule6BbiAUX1qkFiHdJWwHmNLklOOOWyp4s+/mWD+Dqb24VYyHIP
7QtZsWkab0j05H32DpULmQYezBVwCbD1NTJlug0l8BHeO1B1xZDbjsd0lACCNaTj
m8dQRAKdyfY5KGLvGJJfrsKFDDJmLizQwZv4jmLrfNXIH1YLaDs8D1QvZrLpEu5u
CG2eRJuvdbpahgmICNPb3zNdo8ihVZubcOO9HFSKkEWGXaUytJPro6yNVQhcBA+u
btHsbMIpp6eT+3c+CUA6bGd5/hHsTohCm/6RvOmEOc+CQ6ZwodApZlkOffOrHyqx
t1uulw00CKJ41kGhTZPrc/TVxwHo5qbPkreOHWfcP8+In07AYguxqvIoAZhccarV
1Cp05bEEU60Mba8L07mY/QmbbXrbambAC4RO+WdsKLfMnGGgruvXBTFwmgbj3G+6
O/pCxSN9QxO7S9HFqG/0djNuV34qK/pdRlLAAsnhAVKk2bpAfVfGr5oIcJQWOtsi
7GCSY3XwiFtAOMtQsNX4moJa7BOVRM5tDxbjKfZk41rcl8PxB8mUSq75HnEavUFu
7R314Gk/+9Et01gIK5QuTDTl5F72N+X4p2RoQqiIa5LhZyZHFRBoB/MbhX9tqEVD
godtGyQg+jOmlkvKUbchGoKLeqhbOAjWUcjGX3IoJK86KIBmdPdIgwCaj7M2JSVh
MCLt4NquomeBpAZ6xIK6Zcfu37Bli6EoT7lZ6GH9wl+qx4QspmezQ34s1OMfDYb1
BNSDIsqIB/orwBQwJal6UPC7iTiDhJ0lIQKEK7KO9UvldHe6vhJ4YPOAjPKzaV+u
yAsYXIT78FKU0L7Cp0IkkR6wNfnlOWgi3P1A09ecXkK3pBxmBVLRXUTo3pPtL0ow
yprZDjvbbEeyHwXy+cbPmW7n3sYwF8jz+Q71rfqEe/41koVJpKmfpi8gawHYg11I
zEOoZHVTd4JAzozzcbRGU5GW4KvX44vg6xZW+3NjlYgmUzWgoXk1BDMumhsnZHPK
X+Nkcpo4Gnd1PcsZ2utozYWHr3OMqG+TyYYtek4nzOO/aP3PrWSkaqvTUpELsGkc
nvzb86/Sl0AnYtGm8yLD1iiQL0od0O4jdJULOvD2JYomG0P5UYXso3FZWr4tfpNA
r1dALFSxsdNicEnVAPXtQZFZwgBCbu57EKHGaTlJhhxLrcC5cmfIdOUCvjGPjk3k
Mh++wCwRFbMR1cfTu8wDO63koFUIvWeOQOhHkduexVaCAWewXEPi2/P1l5yMWn5g
sX2ksDJbQ381HE9/Y2kRewROYN0cYdMsPJXFqT1lCXH9XzsXAACE7C/cM0c7d8GV
cGZGPacKqoh3INgc9qXzTtR9W/73OSFeI0rJfDgHneaFr3auOHvxotnhO8ARSklj
9ns7lO/tw/CdfmKCaoidnVf6dJaCP5OHom0pfQpD0IrV1if0hYNHKRsHFQvZmBMG
zaxLmIC3Cb43ens7UUXfh0PIp3U5c5FuY35ovOLzYoPVRj2ec0IEsKLRRWSqC/h4
wp42L8/aiO78R44JjLnSx3JtiElgs2i1esGCJfFx1cRMm0ATQluq4MBsMP4wWgjk
rrVIn2zZ9BkBfXazu8BvNnN0nrmXTf2qp+kALeNNeGpCtUaLnOXstBx5btwPc+Gx
qI6z+jg0WHipf56899qH1bNe78MVswMFyjxY0A2iwisbChbDLbHe1Aq/5HsUnQl4
D8rYAJrppn5Px8gKZcE9H7Fu9wEQ0W/pxD2OwJhMbfgUMaipnW4yC/P4P+waHacH
Mnvw4lKqVNLuvaurjYgl31XMRZtsT5UJWc6l17hhidPK+T+dEsYHxwBQmjYMZuNe
OxUwKJ8xbw5gmyFQXChxw5STdBISz1IBIe038QHDxTDWkpXrXnSwuxTaq+enLQAN
tFMqRt7dF7SeU64exD3xbr1WFwZDTbU04gMzdjMElq4i1/SEMqLv4/XI/dZSlAfc
3zPRnbPCexHRstNxMoWmg5pkOp5Fc22VwDIQVX+meel1xfz9BsRa966i5DvDZd+L
OsT8EKA9Ms+Dk+1GNAlvVHTjY/03+UfDQJKD0Y415QsvmBCZwp+ikMKLsDvWV4+R
z8iLjG7JCgORcZr8WhRvaSJmDwh09Dw5Wah2UP9V0LKs+YthimRv1m6zYlRedEC6
CM64JqqABh6cilFiJ9/tcDWhp6sOlmwnlYdeXXWgLYsn5b+mlwr131lJd2s3s5Af
At/kgR8wA1nOluQ+Z21f4LgigSQFyeIEKbg1umU+jDniu0nscN99v0Q6C/fZOjwg
qz72wwOgtcIgvNqdL/N3Ku3SAce370kvXoOoq6owrFh/CoLb1IEpX8h8SQjJiMI6
Cs9aS7SjvM0BaA0MG2vplWLZoXP0t9IFxCsaAymM2qE3vIbWPi4sx0IgpyxORAhI
wo51/uJNF4G80a+kJv52IWg9oj3eufQJzYcuQ4Cbg3jdfKC1BASRnQIvu4CtRc0b
UXIW1YVIAo8DjPitoP4B84KzRGiN8tcBvlW3yxfZB7nufZdoELZj/nnQtVeWQTWj
JqYQ+CGMWxFV18ZOkURloJcqMnURP28sN1jzhu6zcaNF8Hp0lBIQSd4cLmgYsGDb
0eqQeCiYSAT/aMH9q1ar2O6BXHHoWP3eLInoL0WlUJQHecaW8m9cxO1Q4SsENwVB
oqfwyw8F2DEPW7oyKEMsCX6q8uFx20l2RwKZQxWE4zOm1YugAKBO5R6rMDdtMkMM
6JlWjivu0Eqj4/ilZWkhXubfXwQm5TSgKhIJ/5YWq554ldpbwMH6BgibjamHSDuN
IPi5WSe7gQAO3gTQO41Xh+IgJpg31WbmhkIOLwe8QvYfBCT1a/a9/0bXKOaV7knY
k8sF/z0/o3sJApF7iqxzEm+HxC/T20XQDO/2OUWWWJkp7xaZBKOz3N063n97kzH9
UQxUz0QIjExc8Jpv+MBIfA2zrjNzQEMIkGooTE84Gx/PjMOo4jSLcXPggjyclxCU
PFvSzV6QbYg8RSvaefu457J+YMhu5CUle6sAGPLEGDvZ6WB8LBuMJvhyiYj9rcdi
fn+FoVGmxx+nZmTOxp+EFq1d6z1SeHWdqY5ewNHaVTT5vscNOgN5BAocu7auDOA+
XYGAWYQGheph0fEh1aq/lDSQ24Br6Kn0cP/ql/OIMYa2/Hrmmn+ByINVoaql2x7K
f5XxGdW7AIGooUJdgVtBy6/jgztlZkxQ1Bg1fP7RNtt+pts/fAzo9gBfCsdlsfHr
cubmxOd9MVUdlLRIyqUo6gTSX4nJeCxZZMS2g8TFsiXnK4PL/tnFRoq2QXL8//2w
vuoQbduy1ol278OyM9sI2EfbWYVyF+6OQCMTDKyoGr5sVJaLAntfn4jwCIUDe59q
mH5uG3mmsnRT1Iwo29+1RE3vJQIlG+wgYk8+dyeDAMIz6y/SznSZpPdZp2AhzI7w
r1K5pnI9OQ/+rBsrp3cTQtKGlRoQoyBc8WGdqi+O+R7pxc4blmuaLlaT49KkOXDE
CM7FRVzf6DZ3JPUcdlC7Ok4DB7RPj4s+MZ+pSTK8q27F6xc1e4DtJG6fVYR7ol2u
K7/Vcz/Z5PYGidFf+v3ZF9K6ZKsAw7SdwFCdizuZMhOPDLkf33P/8bvwI+nrRDna
W9cSXqKFdIUNKNjHIA16KwKe6IgOBoWczIhobFbNih7FvseoChCnPjK0fgHZ4MIZ
mFA5s/Kw14INCqrIZ0dvBH+9chVhYLCVZ0oS5UmjJd3AbRrlM2hgMScjyGiZW+Yi
XnQtASJJG63yGpByhb3tDrOT1KeIOHbuNFHIOtnAEcjt3rWmB3Y9gwrewiFx0XLQ
vLjT9ysqt/FVFPH6k0d8ca0sp65dMJ1Jm4qndEhUZGWDijn6bsRb8IIGpAsSfGAO
+SZbCT2hANfSqEnMWleM5ZCValKu3jyFjz8cSv90FHkMvwxoZ1iw2knM630kf+qj
lOdAcWQJlH2FUmB/U6amZz2iFsp6iADDjYU/VfDCqMvL6QYRi2bj5VpNkVjduXnh
OUDlv+iNCECHCtgi/x27+Q79dlqAnq1H5GdL7erIMmjjl1vqLxLKsyNJTgqWpFot
btj8+OGT9LVdlkveSt1iTGD5O8thBk9c6X5+aBSrltJxOcmNnp/kM4o5PoS1qVDb
8Palxpa9JJjmNCd86z10IQGFXH/dB94dVctM1Pl+HRW+uYOthwCdk0pWO0aiAc7u
iGdx6y21BnvFdzzqJwz6crPx7Zr1LTuYLogzo2PSfmen4PQKzJVgEMoh5Lhg5I5f
ig96L/P/3ZBVJ4QnGKbQn8hO2z4pltqCoFMxjYFQgqAARjbdWtxNTdMEn3gvl75x
0XBvHsjfqU1PPOZ029TOCxzOgZrydp3pK795nKw4hHewnWqEg10HqUKUoyMHcMCh
BfskqyEuMYtQI/vg/ZWV6gx/RrxE0w+5lKSDXLCMImQStmMuitYTLb5xKJ8AWsHE
8BA/oVmOc5ShkAq7ng2jujkMHMj8st+0vsX70Bt4Eu6PpStVttHQRRABXd7/Csw7
fll7FJjkE+NzYT94WGUYSzFdsFQBK1gn7VIcp9dRBIdYU9+/jf+39pItS6TEh+qK
Ktb8gvILHyPU3414NaDgpo8C6bG7uJKz7f5WoX8JNSOt6mkKe6alpD6GJtsMSvQl
MVIFSuVH8D4f8LEU1DflAPP3dfEndH2CQN9ButjLsT7LZk9F5uNYVDYSiTI6DTXL
n35fyECUf7iRM+S1GKoUAWCtMWuUHDkDAHVpXRrRxMseyiLHXNqPr108IGZenOrq
aXhVqSJL9cFQeiR1v9UBV2r7dB/82NcxfyUYTW5ziTI7xcvnsKdvDmkg5VD3RkaY
wDZkFFB367YlnLJmqiRYQPiAOmGAZ4R9fJ0v9NWgi8ljkSA6Bqwhqex53Sl/W6fP
GRJBHdsOJUQkY/3NEyr7UWm8G8wvl/GS1O0QOsSLZIAgKl8323VXtiwRRluNghY5
nuP+t1nj1OfkvwjR84p1ExjZ5/bztZ8CYoc31uSdQ2xYsJ8y2MC30I0CXlW1pduZ
czqTLjo/jfj44Z00HKmWS+z21ELvZK0byOww2jhC0VOh6QZBgAOJqtgKVF5UtodX
rL8+Nyjq3nso3u27WZ8U4EDqZaTCW9K93Hd9A9drdlx9dAdFYnVjUUQB0TQiW+Ro
AfO8Kz3vspiH41KRfblOD8xca9pRXN88wwcQqESIb4akvrnreUk11jxWW9bnSkmy
q1vxzNCPaQ7f7whF1pQ1BmnCuvfmWiRSAOFKAmZZB2O+DWWm33bvz0aNW99HIIrU
o40i0JpHljShZ3v/0dNCTQQEZFj8mMRa5w21Fp6H12WSszMu39rmnEDzY1aFmKq/
+A6ffQ6Bl1ogqFuRlepGkSvUXcjcQoO+ClmMchE34nNQ6Ax0NHmdxIqYIcDjnQLI
MY+XTX/cAgThQlibmSlmVy/WtH4ha+RufHwsHvgUg/huaFJ4iLITcymcG4VeDO/0
EtF+i7zPmRrVNQQNkitau23/hIR9r1tm1Y2MfE/aqg5fQO3upafePZn8KuwgbOc/
OFJz3kMCGWGWNM35vrY/m2ZRphSY4pKxQA+p0q83lcluq4TKntysPSJyVdluaW9S
8iD/ruwkHLUUzbJKVreUUR20SiITUKdOGtjMcQ79x0GgsT9qjbUXSjMBoLR2Uht/
AsNlSKXshAV1N7xsFj2u7VH1HH/aJh/8zGvHn/yXbsIeUQjWjnnFdTPW0ePrDhzb
MsDg7ZniMqPS1+B5wQv1W+BraEpev98RGvGbqRJj+ieDZawkGF5U9AphHGjwnONP
FbJQuzmlZRYmIOEVjr0zXVSsR3S0v+U9DDpwL37PbExScPgaEiAhyb+tzinF/rff
C30ZCnB6hJ38ZCJ4IkoA0HW/UiHXuT6SWt+F3oqFv5mJ/R/I9eP14RiUgPK/f1D0
LgPaaYWGBoe/p9sQzlEwMxeKq1W+kmyAiPMhPzKDlxVDWquAgRsCdiB51rb319lV
uhUaPjARIpnqyi1Dv6kzzGNj4jvvPO2COy6cB36H6MFIbD1MMDn+WOKYMxCwdAjT
ArBRR6FLpsLeNd7ZVX1gsuiT7O0W4JuUd6nbFnpfw5sDVbxguGV9UNKIVy1INmAK
5bDYZdCovnL9eVPs3lclFzKeuXbGpEagCVkIj3ngTz1+FrMumOtKM2b4J87+Fs5m
Nhe0a7B0rZNMvQTAboYMFg+3L9oF1M8V0CjDGPTimVaBXF1m7xXjluviYrmzdg3Y
MpIyUgqG44OD7oHgvmXfPkh8qDx1rhZaF4YZ1vEi1gSkP1Hh0Z0alXtxDDhT5q94
bWynTKLFEuZ88Z7kmX4+d2mile5LcmiZECAr6ZhQMRxC0iCEagPck+pmUrlEpllC
3SdxZhta9qcGK/mYwC9QnTFn9tkmFkvVAPFeyNCQkb/2UuZ5CZ6c9Naf0tpV7zzM
R8xMDiXZfEOqgRqDjzdvIOPBxy3aMGJzPytMjMfrnxsKO5zvcFqgldeH7bl3AuSZ
izL5nkWQjWWBl5pIes/PppuTUyOcABmvHt8eOwsLVyuc7w822Am0M3cn8mJ5xquk
XYqqGzxNRxeiaDGhSVkjFo32T6gEmsQaRE5BQitHkcOTKWw4Y1hhl/v9d0bgS7vv
JiIycmnSSBqkpakMVNmfCJAjpwTx0N43u1Mv1pfF8WZOzW7xmGnQZZFoOOtvYMax
n0+xPon9walbY/y9N/Z7+70AuH0wE2xlMMfn3JyUNEy+ipuvQiCH/SN5mK5suOhF
j15JVWfjRoOOrEdtWGT10dP1nRT/cu8x1i8Jred73IibdDTj23EIs2n96Lp1/t8V
wf/q6UYN9pMgsrhEL6vn/OBDDPSTKv/kpduWT7telfhDwQcfNMEltvSe1Evya1HG
AZfumNqN4uUfn4T2M+H8dlUyrDf3ZbzCbDjOYrZ3q0IJACtUDqFN638l3yD9f9lI
g2v/A8zxqww4fuFAQBQ0oWQwOIm+VFCfwESOHlrNHcwjb+b02ZYkKOUHgbkvaObe
q5UwIa6Z3qIXIJ840dmbNlnCTl4HZAJf6IR/XgPt5ewbj87o1dKfjO1cv+Y9VDxM
oxyh4OMoPc7rZIi74fJjIgC8byq/msEuhaEekJnGSJEPIddLVuqp9Zs5jaqYLXxU
ktUqagmaiR6nIwMaRmNVgqY9ISmFB64m8XrXmnF1BLRUjAb/xdpENfQaRejmMb2n
/xQmqfZvjnngFEwGo9rvW5R5+jwggvA7fphgHnsF117K45NjtH+hu4KibclcuKr1
eAGlU6ZtQmR55eAYqdLQ/rsid6VC4wj3IsLAVkdR1pgTy1PW6zebhqDxZhMImFdS
vMQK+BPoPlds5i6opC8keyjARqm0tdHtuqjn3g82gbye3gX0OkTxpoGcRKrBIoYZ
10xBEK1TQb8g2bKHnExrEzphBCtkxc7epoUrdFNCucIiGQ/pIJeBYYqabrbi8uaK
AxB0ig9WG4ooGwzjNqEVLDE1zRLmvlskmPma40zwjUd5ArrzIJPO8aaOQAL9yD+J
dBmZ79aG4kuasT0j2k+S14GrA7qSU5Pg66y4PTHDpHfdLzQh0XuDfHCD/TcCpEsz
lkI22lhLuJ+GmfUYC4OSGqiILpFuFhJl2H483E3fgHCXbEx1lO72jFe7d/6X9iyR
BDcUeE6Dw61SqxKGYsf9WPBd8Yy4YP6kIrUU5c5MRWOlkTODkLlHdmtu8VImftFT
xuHCPR8qirktyhnaHe4avK/RPOEunxuJJWxlieYFn31Y1ZuJ8ylHryBaU55MudFO
dVOXY0Ud9Z8te69SNcLtaoSKrvP8I5NlrekX+QP/q+la1boSNAY4icBGyy+2SR98
/oIt1ERzid/1SwhsBKo7fXl8+o1cGsLO8nUDUUfiz8pEP9RGpoVt+CmY/Uuwjedy
u1Eu5ah7v7wQM8fFhyWsyFt23BGL53GQcHdnRFynrZi55oTmAGWALN5dQmVNUCzf
JW67ZL1noNMMKFauzO1AFhq1drgAwY7Azf6JSopiSfC0te8iK5q17Dqk3SD0lFKR
bGse5NKukQ5Qga66Yz9t+YPp0LWvmwiGkm0+sWK6IJA//OD/HoDzWXys3dJpeJnJ
e4cHNudwDJOb4iYU5I3GPsjD7vNXNllqwivUyoByYMD7LiO/WzO6Y/vfZFbsHBA9
t4yVQDuvGP3rM/JL5ChyhpqAumcHh5hfuRpMlB1ZOkuP5nsBOGD37AqAhsAvQzbn
yFJtodGYv7RVjRvO8IBe1mjoSJi+fmQWlCyKFPIhKiEu2SVLU8Sa7BtC7/AtJ1SP
s8FtE4xBDlqTfCWHHCh2lS4fbjTkNGTF+rsuMwzbmkbOwkTDJkRbybRxrGvQR/lE
75RqlAJFiy/makTEHZl1BPIwuK8dS2DmZrJo6GfheA1Q0bRPeC56x+rR1e8lJVOF
OWR7Tf5MZnEBL3KQoBaIvH1rwoYmLRSJcZk7kJw/lsypiH0hEQ6Epr/DDAfgqfbN
bwofGLBVfg2GS+uJ95Kg7YoMu8QZ24iUYvSaafx56zQMXBMLy/fp3BC3c3CbWO8f
Z2Z5RZkZBX1xKydswzhKP2bGq78wyR+UToYnw2G6l7UizSeZqhoQlQBC53DKvlGH
PdBdnrnYnOkLa2wiT/JzxX8wWH24Y8VK3fcdSD300+VKEQCadGns5uGQLq8SzHxZ
PkQK9xHTIs/xuJtEFcoSdLtsm4IJMmaN9nQRdfvGPAqiK8IltPQS+ZxyXri8dY32
eXY2toq5WhVRKQcjEmSw50/+0kWE/5iANSQLrh370SmhV7xOY/XkRxyIZn8t3wJP
+0J5NoA5iOFED6YevV8TBwS0xIGzUA5Vh4yQXnwCDxXFn1N99eh390FZ/GBmdmjL
yOFSIXVMXyKNmJMI5C5R5zDlz1scDdRyoZbvIChqzM5BXPQgFDgcZfdSaMylq5Fd
ometzwEQOayBl4zeQxkFhhI+xMe7ITK1HzhePfcXl+U+poObzX/82wz3C6FKkaN6
YryMU8yMADLYtpg0GP2UUGqt+O5/cjKhNP3MIBqe6f/v6Gf75+Lt8M2r40D1ozOG
tWEGgHk/nYt7ToFKOFVaOeK1ikiXNEX4/PudVaTUS/biYKlq4mqxS6qcSR+NvlgE
NPFvURPsgwAyzwz6r1w2jkjujGuTPIjLTVFdfHqN7zXvqytKOjhv4XOqrP+QCmtz
cYWiiyDVFEE9st7y64T6vfG38hpaq3XSjWEHnQVlHaFsrMHWHDR4zeBsLqKUakQI
Qr9CB4mSozB8r9m08N9I3JuTaMrtCZGQ36CLqPjSXHziUJHtvzT7BuolD5sVJNPp
LYiMl4JglCSig1+rXtiyBUacKgY4+Gxa677akbMLpZeYRRwRBs0Mj5ADKw4s8VUg
Xggj60GgaeCkg3XsMnVQnRWbwtl/6p5Ej945gwogGb8Lj/53d5uwm5hSUwCwndbZ
uSSbDFdgmmudCOhrKy/XHqN1D/FiCdYLJ6lCF1ekFW7gSWzJDBuIMNzQlBVC29Dw
Wt43MvquJutLATQuHLERNFu0EZGZExpS6e7aPEAM7uDGLrdgjCc+j//abk26Jvvm
Ri3sj/yEHdvSz0eS0ne191CIU/6qFQzkhRpzCvISqvcWrxCi//jeSD7VZV4RkfCK
0UPbIHqBdh+FW3Cm3HbsZB66ls7v7If9DiNYm4wzXZvpvBI3yp6wHfKdyrPkg9Q6
Q0QdhgP/tX7NrKBNmNwuKUnNOptNqTAGcvoYG/8afPc9bceaR9WPvcyV0aqfriHl
WGl5VtH72AJvNR762Ax7ozuCBMiwNgJCCt3iMIrUEdJd6WMKXbapKuAQfticEdXP
2IOiOq87awaFyQgZeoqxRHk8x1qfJeO1pFd+9JY9pYK4dQ0P4FHSP4y6zNb1OKwu
qgX5vbbia+AOfyyuU/bk8UAI3PtRzZlm4hE5gCt35LfNzUgUDTg8qTfkpnPTHZlf
tfO0k3opBwjeWItNDwcLQXzHW34Z3367RM0cwK6B1uAngVlpiSJC1EDGvxXM0v+P
JUHjl/Ph2yVWwnJODfhl6F8O+rp+zbbsgt7ql5ZzUczuNhHkOCFAj1AzRzHvNrZ4
YnHradkI1mhIPAOmdByBlFVEzwOq4jSvjqyLVTwZhZ23L40ccANeOANvqdRI+v5T
Ag2oBjBIVYNpdBkhu12zQ8YGh3JgKO5QYhnBd243nCVj/3rbd5cI8o9krnHFJd23
u/yfYCHXLhV7men/i+TZmZlYjOsPVg70XWYkTtJrm2pMIwhAvHvWvjaRIYIV/bq1
zo0PK8rm4eYjC5iG2bYd0zAO+Vr5rel67jJZZ3HxCehtykI9ZrO+dL/P0ZZ8VFKz
h9fJfmzOlovImqCfWCio0Fb44hpmiOcKUIzSKdfSic8YmnbwGm3JANyxwOBk9ciW
wGLmyW2w1fxrBxKbNhflr+6wahqBHRD7RLKiepdgbUhrlX6Vs9tgCHKce0SsSflx
D0s/6ph8WlONZf4M4OybGaX1/YaSTtrnHsNaDe9i1cUlF//ErY03MC0/gdlSS5ts
lC7QrUa2vuWFrFVYtYi6lQ7TYPZC7LopS7qTH5hR0II8BFMLx10bdrUgAis94eZF
9n7Bv3s7C1JajOFHTv0BlEl9zOfqazWEB14eu4VST3sBh4m1pdukl+v5I/nWXxt/
GadekgfkVhA/j8hyofdbzOwzvNaeMCI/H70/7oxy6ud1BQ1+dPYgey4d+yZIIEn7
anTs/c1rEX6tO7JhJ7LXHR2llmlA9zrpojtqG4MWTaSFUlxzCh84Q8NyQHtqYXzX
tITVC8kqqiAU53w6qBTafOzBtYvOU+sPZ68Mr0kPPBDcQM7GODH92tVgU1+pcFRX
W9glJfxAKW8jc/BN2zcJOoLKjx2GwxLLrQKhL6jHVWdRC+VOny0GAO+cnBGStETo
AHmBKP7zdkQYfcTBNDrFPhEq8MNtvQSZ2z6GNv4y2hEO48N09se9U0MnYbXjkt28
DPZAENlakujm+PJku41DPnbkt1FnlMIgxpSqqz761v2x6Yr04hF0i42Fq1Xv9dtp
L2vjmeluzNGoT21UYuNCnpp42DCXqjH+l2wM1Hmf/U68LU5kg+WEzptIIbqm1yeQ
HshFFC7zgcczABVHoAw9SUi8S7NTHv/i5LJ41qgAHJguqCf46StoHAgAcUpiFnh7
TqThRUen4eJHiC/V+rfkjbkI5LhdAsZlEcuX/0AcSplUXAjr1SceXIlyCe9uR1R/
POt3tcmcrJkZ4vrwDRkBTw1CQkvMTwU+tgab2h1k+8Vh6VYe17Xp3EfL9USOrjgP
N0lJcglnU0KSuy1PasAsELhRAbyQnaWk/lZ6+lPnp7Cu7zoPclW8V4FZ7m2tV7+r
S4QXd/gKXPqtfpwRQtWkcMX12hhOLGftWU6tr56XOoGXoF0REOaSGut+Oy0ptBZn
xNVy9OAS637dYFI77tx5bvw13jRl72zOny57FApugGcdv7BpaCZJ0W9Oukp74yKF
y6TBmxCzUwKgPciG9BJrWi3YagijNu1CLbDmcTo9JwjIR+bi3dNQsYA8itD1x1dO
R70GcJsitQZ4tjv/kErqtk5ROottS5vCiyjmAWtUuG1rqJrGG1ZvwI+2mI4jLvlS
Nq1x6mBawFTIU6klA5qN0uprNHK42erPpTh9GzVVEeLCRYPelYKVaonVL1Qv2tA1
1tK2oA1D7tH09IK60Q86bO7IM0ArWlVVUcfb1xzo6rmsCicJBE/7cwoQdn+qXoXI
kQNTroF2ZslmL8JTxUGGQkwPvAtCPb8EC5Ix8gDyMA7ZkvhkWJRqpbm2HYqOdFf7
ec7fo94AthI+XSdF/JwXAYovbbEgvIrCY4kVYmw+yui6BRmo8NtljY6rZvjiskN3
T43EW26cBFiN5ferNclbHyP6JqL3mOf05ZFq5oH9LluULTC7vvDTOwqYVKzWp+iD
xGqtjofzROPrKrSjXNV76FjWm1MdGX1VcqfW5VwLwBNO+R0uRg6IFlxDG9Mlj5qi
Ot/u6AixT1YQuo3zOohrOhEKkFCXatKr+3S7rnOwYc9+N3RVc6bvqb4q2doGVsXU
Gb/LQJP+GRy7WZQQyM5qsgr5fdNccuu+lxIo7h1tarsrBdPcQo0y9hAeUMcoA9bx
7bKi3ov0NtUMfVfW4oibWmJhkogSmh0VY85li0gu//R8zAS0ofhlg4lfYutWDm/j
NEOe4gjMbzTomx9EMAb2/5OBwCbmpk+5GPsVIVQ4iqSoWSwmXxjBljF/quptsxlx
oHNU24XlAXCOYu49EXWRKWs/y+sotLiqCXtO5FdEkIYo5fHwdLC+f+oW8+jCr11b
NF+7IsKxwcbpNv1sS9aken3OBNBofC7OYBo7GbSqg3FoS8jDswCaygor3kUv3X0i
5uWTVpSz5QQvvC9k5SUIDv0R/Do61HtfdaUu3BbwJYF1HgCfICcGrkDH6Q1/Yo8M
BOaQA+MZw9svywBK/LUYAYHXOfGJfAuaCgOiMlesyog/xDFpE/pIE9jCXFXboj+Q
LnzC11nH24jOhUMFmrLAGuWW4FnGK+Cp3CEDWfnBxfQlNkfc4Fcy9bZ2YvEyRCVC
401zta6+qlB+AiTC+VdcHkI/ro2qwlnC/JQcJjITW8tol/t2N3QVYRIZ/TzhS9P5
cWUR3mxFuMOD7wo29CrMqdGxfbZZnOnYIo5xuabQQeT+urQrxmDyFWZV9Rxcp7Fn
mMOh9Bmb48ODqL4/012WX5icEdjOQbjKQh40+0f3BOen03KPwQkOEXmdOTR/haNa
Ph06HOsKIfAOAO0bEBseOQKz9CnHCPpn6rO92X2jmRGOReXrLeiM8H9GqQOf8a8k
UQ/wcy0wz+xbIngw8XlSbMcJGaxhNQGVLk3afsERSzxXN9hpiKkL8yyFD9bztwbm
r3Spvwl2NTi3XTYG8qlVKsxOBJ1+1LSxzIDihLhutPr9JxY15bUsZOKZMRrGDX8z
vY4U/yMfszBL5GlLLxDksR0ihX0kUZgMq/oBRmARVWqh9dl36jgRKlZHXXGWlalC
SHjflY32Uac2M1OCeox2gDiaao35cQ5nUO15ZRr/nspUuZAK8YO9tCV6QtTHVXg0
djoMyQXhcLzK1bsRgyzJAYvvJBnoK5EJdvJrQpMnnheaZd7S550GPK06i7yRbi2r
PzWJ/MvOyGZDWhJDVXFakN128rUZeRw7QfH7GqdwQ4E1AMnLou21HA+TWBF6RjEb
NxvKNnyoDdACeqxMG3O7UDS384ypAUxK4QZhIrzWLumhpVw9DtPsyCGVidGTfcxp
4f0yo0zDInrwnxwqkBOvTs+ncrrncsV8LXrto1cCTSOzVrLB7cfwAwIRBZWMiUm6
L6d74W/6gPSdDUKQ5qPpkt3y/IYiY926DxeZtBGG8aZhvgLQUjV0XUlSv83aY0hX
u5HakiBXXDW7LeZef5E8lNe5V84t3TPYCniX9O8IClZLNNGWCpHA31e05TNs5hJk
Xae5x+LKutQOol2ceujNx/rHamou9/4zoLA6BJSGLKnw3ut2+oC4USpIFJdQaPUN
LH4+21dOJ2UklHQc8Hb9fMeUYkPeTtcbLwgJGPmPv3dlBP9wl/Ji442uuhp3JW3x
rwEt/e2miJYUMLLiowr6Qhs+Q4JtYWPPHyWb1tTclLLYv/o0uBrbYyARyapNji9d
yaPMDZQWGlZyZYCGPFj/6WobC6YHyJkyC4mAnpb07sc/vXdS/YPb4vxRqAEUkSpb
AgWIUpfPKnqGE5R5BPbsE/M0768IF87yKH3g3E687nTWX7Gztb71gPrukNg3YHd8
B8Av7Bx3EwFy4LDZlsgiF9DHNv94IS/hP5PfmFB/WbZ7hD+6pUhXGGe/CWBQIGyF
LS69FMglawXN1nC00MVR9qN3cZ9LgA2vElWt0KKvvDCvnynXBOL6p7wTEqcPVlqd
AOYOQZH0afg2bP8mtuo+IIrCMO6JPyBLH5udyYet84l+mlUG0SU+cOFlBTbQRpM2
0znKmXpMtTVdpxum3SZpcUDXi9QTqjJVlmdKNo57HnsIsuZIUqTzY+MALLG5h00S
szUIcWlv7zyDnrPqKMT4czy9aRUQMOQHvQpzLDcVXHeEIM6AvwCIJ7XcS7ilx4YT
2lP9emfltVCWEnawN1w4V0NyiTi8W/StTH6Zeze+anS4VJUoARI8sjBFnZoxir46
EU50Nf0MYrjTtHnCiq5T6TXlchrJLPV2mzUGKV2B4nQgVfBPQmwPLihOIgZdoAW1
BmV/zqCqkO/6Mfl9N2Ek4ydHslkzU4tr9WeIYvfzyQV2AZQsXUKX04xvVCluOVvm
3ivKzu3It4alZZuQLywgAbRpXZSM8e9nPlei1uqTjQIzH8eCG56QltFwdE3Oe0p9
+Cg8BoBjdkMzhziC2UfOmAtX2iwF4+stJi6/b2UbQkZIqObnD+cDPtKosiPCwXIa
oJJz2+lcC5Qke4nlcXIbtcGGZ+9lhxzewcJjPXWUtnrmR+YTz9rCCUgzh947G77e
NSQ9gU8howL/Ab4Ev7CJS/ovf956mU1ZKN9r3g9iQ1ga5O9X130DSR8eh3jkKFMa
tt6v8kFIUNXEZOV+qmJeeVctUR/OL2/KRhiP06F1UcoN/xTd5fMoDG+lm+X2BIp8
7DScMhoPZl3ThOf5VELp03xgTx10fYmWxUCaoHF7tEA67x9DUlwqimK1KbbFZtWY
N3p8aQRX+li86KQVY1PUGQvIuqESSDgHmLoOAPQjb+pMrgc576GuWgoor5zAYwgE
4M/9ebjjhis/aVQxP7Rgm+IqdtzvRX6BmOK7EWd2P0C4Vz7vpkIpqBMDRa/5OJI3
+rhZfmpWmWZwsKfqXUt7I9EFNg5nN0unMZ+Dqz9RiJJaJGccYDppafcSvYxDOeiB
6HrIGiBgLvGwTmy6k99+7NVv7cLqJT5lJGybIfFObAwi+Tiz+osJ3xu/uxp0L34e
uWFsw2r4NQSYOGDhCq8fEvPe1cV7wmRXElbKYEPDQhdk23BA0EPv9wZssX5l6Gk2
+WIFEvXqdF8NZ8tDZUMl+IY9wwAW3cpjgRfuXyg+fuymObvMwdRoySXkstgx0Nug
aIxPfZDD4ktayW36JXqLj/WPOYutOW70srJxMpKCSX4dSNFhTMjf7HQh/tCWfXle
B343Ug37NCvfH6It9f3dfgEEDkQyC+swQAKnZ4OP2T6zK+s1RyOnl/MvsmSKxyPP
UR/ZoDdECAdxuimf+Q8OnFEuhphjqMJ+ymP8BZfniAKPX+WXgct3WaLXwsIG380N
Va575ympgBlHsKTGs1f+rmZ+qmdQKQAYkepPXGX7+5gpq9YjLOpbPmKxPgp5GBbN
WBgpaT5zF2yFa9hwF3Jt2nvJLVubZqgtBb58/+JRtlWUh3TQ7VkOgui2t99i+gxH
GASBndVwMiq6WdGwuO7LrQPuFMwo4u/pSM2UxuW76+St4dYhDZBv5usGH7wT3QU3
HhuNTSeDB+FLdozQiBxMVEkLaxTeORoMsbBLGGxtW2FtfzL8Y4ZnZNK9RjOs8T4D
AaqMbHoCObhA9YCMqZxwPQmi2Te9lvkRDMO9Ju7k9vr9upT4wIxkCrmSIVzPjwzk
QmKmR/yIOtHx4bQbZ+KUQVNGgLdf7MR3++2ruaMHj9rDLKD0VrClv1hgDehk+8fT
mpAr5GCX31ZnxNsZAlTTTQP/DcFsv4h3tMXbe0CpeXLNAlL0NhA+0XsM9nWoTG8V
IaKIdx4j60QgFL1qHmn3PJV8q/b+h2lC9Mhg37YsiTla9uW5ampiaX783aj0M3/n
P1JRHV+HQIwUTksLpQvq7xKJ0bFFfUUoP3NALzVox2L5mm8CQHQV+TlrYAj2UV0c
5PcmAE+viD9AATAWd1KPkB38rwAIl/3FKA/Vb9YqGdL77g2jUF1/zXLgKPqPizJ6
arnPEYli1DtQ771mheg05tx9/hGy+ymb/u3F5sZwElmz1FfBz8H4GKneNzlz6+qk
3M7MYu5X76HXbvRQPd3YhdQnzaubufGJKvR1DIz9BYyt9AuAxiRjo9NWhYDIC9Eb
7bBSmoP65QFcYpMc8SL3FQXxgOcHlqACGuLwCwJIkX4DdGPcJXeCvGv4dqIFqWny
GYLVqBvpBFs2zchm5Scjr3W7lZWirWTWL1SAtgi/k7MVMOnBZnAw3/6pIKalUu4w
NHJxT1V5zUt+reQRCzoskx81uTuKVH1bBIPbGoQHmGc/JRm/VqS/Hxe6LqV+mKTP
Xq5qavVSLakf+kuuOk3gELr8pht3xg5MhiibUI1iKNj0E78A6BJW8DWZfc8h6I+L
PfCBQFt+BC4dNt/czo0APtlzqX63j4dVQEd0gtdZY5uhYrSn9ejZNJbsg6fjlL0P
h++lgVjD+BEXhkBXeMLXauoy9/y/lxanPj6SlHHVxWjx2wrNhDlJ8ZbvldN8w+ih
bkbyKqbuzDEqSHmuOgkscTcf0ukLECBa36zqbwTufbaMsNLG0BjBy7KAjsBCbriq
D4EGOKv/tiCuFeNQM0/rWoL8p62L8+vPZrIqC3ycS5tOH4q5G/64HqsB2EgFDr5z
ABVh1GSNpZ437Pql/6E4h2NUu1MUhDCx41dTxM97tI5zVqQFgV1sohFpTJnSJJ3c
QRvXwSkZVd+WbKuEh6bVw265mypdTmNqYxt1NCeqMCageVD3bUzckVNEDF7rXwM6
buMf8/yqtsUpwCMONerYz1z8313RAUwTTKREpgpSjeAoPB2PI2BlmpwuKPiWEF73
1LUuM0o2GbBmJJMVVxmA+WdAkJBzDLFVlCzo0rWFAWgp6zTQCC39bQ7fiiNd5+8t
w6HWB+a3i2Mvr43c7r92eckL7E7felqFkXsOhETuzcMXUfER6l1CB9NQFb+ik0k2
TQpSX/r+ko+Yy3jvh2U/474QqdVT+NxvlC125ehnZ/aWvPG2af+2jZUbVKsUvZrl
kUMjsUIMGVl6+TY5sdiBTIsrQimnVhzRUes8NBap5jHb6J3FDveE4433BF+VVueA
2/VRvxYZOPX5LwUd10MtWl5dtHw6Mr4xJ6Ob0RdI5gBqJqWxTx4+/BTup4+mcOTM
JyefALJoM6obJOYdJYs7l+cYdqZ1YYX598ycvMfjDTsXlx+2lI37lUyzsEDZu+te
rOYVc0FYmqdvR3iDRuRGZBJnnFtq1bLdo0TazKUq8MGb7ZMBQK+EiUgVwsY3EB8R
R+ONSLH2cJoyiJgXDUH/t//FfvtifVpXy0a04n5Ifs9pu3rAc2lcVlnjfZOKNh0a
EpJfM8cySSrJh2R5wTISq4E+Balfo+HlmNlrvVAdv4Tyy/up35XQavx6vDV2ULyf
ZuD+t/71rl/o/xBwSG/FR8HbLmtQM7dcLHWLM+fhRDd+KVb5yBzytx1s2Ul8EMZf
ijFyWi3MuUMTXwFU042f4g8vb5uEQRqpZwn1/CQPREJ1YROrSE5EXg2RCXsfjNU2
rSCMDrShxca6Fqdn2PJFhVcS7DvFAW3oZ1cceys8aJ8t2xvlQpaBMC5ONrMll1B4
kxG8TEkgoKTy+uzm3MEzWJM9OpW2NKkuIGdCUQDeZQsW4BV2IAv5uuzUqFqvMkXO
M7iiRd/gU2AZYWE4qApSv2ci4MFvwR5evsTvcfoxTae244PdQNqVe4kvYKt3joaJ
oMZM0ML+HAB82lKdZSuXAwkM95jILM51sdHgn888WMS1qFeZRSVmrGcFjWlyQdZV
h6B0KCclV31LyeFPA32Lb9iDTMfsgN5tVsMv3mcpLuur/Q5XEqw/sAK3f24fpbDP
TGGFzpq8tNqaafeHW/HWIISPaT4jnf9AzR1qxnU9nrUeKSVW6cEdikLI8BHllWL/
QNsW2dQ1nR8+saBigddouOx/LeFMIpYkNqjatJK9b4MYXrP284VimHXtMeKppnY0
aT6H+8h2gsvgINLhu2YWA8Zm42ytYeby7XEPOIlUfadx2G0JiFHAKzJbZTjVPEJV
aMp4W7FUryINZbLmsPAErStbCfaUUhhxobYbzqtxrlFPnWM0TBVsNxEMowZS2bEi
fM+PNeyIiSZzHTl45VTOcjvEY8wkremLHbSDO08g94ieesAaJfjkpXYjRYfjKTkJ
LWT7w7WKwpKEral9v15f5H6qy5VpwG4Zql+wVZvrMWYXJJ88Ad32H3rObRamnLcF
6Twm8oGQVGw1xoNeDyAxFMMu5vkleJuzNJ3vHUqPTxA6vzAFqy4a5OcXhRUEyFbr
nbTeE2XrK+uhSmoB7Nwp1lRevh2k9aQP8vRtFk1Eq3SydcvuGrFitoP7QjvBKmr4
vjksLnfQashfUuGDhyKVUjjYsJFqQ9zPz+9XScThyJt/b5TbrPPHr0GCYtSr4UwT
vLFdOoTvan2brFPBQtF5RZCZ7BR/KkY2327x/zbjqSEnVe+BlPu+eMEUuC03mZof
Wy5iq+hFOtUDwjaQWt/xi9Ob6W30493zOyXp6Rj+EBUzAc2P2IDwuCkhVqai2E5n
8W0fv0Y6pFCrC/a5HpAemLrQLUEe6qmjJ4HpJUn2gOnKK8bD7yWKR0yoSGYk8oMp
TgyvXQudKxlcSeQ/W+Opviies2KZWXBcMWCgBpVUJOUw/HQ8QjFphxysNOiq+zjv
tI/FBBvs0AX6oOIVw1DsMBZWGk7CcQPRI+XB0aLJuQoRBw7OxoxBh0tpUAQlvEyx
NJ3JCu+jSfBj2Fm/87kzHOONcSInv7p2FvatAaXoZPJQhtLP8/d5O/NjRTAZSUG+
EG2uTExCeqndSR+PRXJdfnJnMqWCWRQeDpZcrUG+kE87zU+MY41WVH3PGX8jBncw
v29ixxMyivRo+jBI0FVZ5FyE1kIKL4h56etEwZgY1PZ/5bdS7rqsjGn1Jq7+awNc
s7ssmfe15FG2ozwNZMZyaY9Sq+srPuW+PwweENjEhUg9NjVkTnoolh1XW0nOzYE6
OnKHH3OhZfoKMkpbXbscqwYyy7qyK3TkAkZjb8l4nKw6PUBY0Cpc3naGHxNIkSzy
O+rvWOdoGpWIU4OL8NnwZhcFFJC4Dq+xInGzQvaiTgyOCKQAhW4+48NDCWau6dXU
wO9HAv7nXchaLiS7+IjD1jqPF0rAVQbeKjp8LnL2rQOEQgNzP0XkUXIdIXd3+aII
0Z+SqZ4wePdAi/J6A3ywoqwRcOfyjivuKdv68i+2LX0GBGgHN1qxYdpb/r0xR+eD
RZlOR6L/hz83tqn4DjYA9OUXoyI2FQeQ/D2wbrT0uQ1/BbsKdqb8Jnya36Vkrf8s
9jl87B7mf3u0e3LeLhO+gLvvTXgTvGGECFQLCsaVxLjonS1/m2bHERdAWlWD+Eib
SF/COdG9KQWHmTEONmtr/a/f8DE7hTo1/5H2KZj6Jmw9fqGR0WP0hEp2riBwtg07
78d/We9nUsPgj0Ul0omdI+1/MgW/EmyRx7nXoapn/itz6QfK/CV4+zh1zxr5fAfC
ueCAhFWcs8Gz0z1lstw28lef2+bx8mp/1R1RShOpRDvVQwRpiy0yy1azvw+VleCD
CXQt75SwL6y/In9mSvVx3sXRvSrsLtPvMQfWxb3NVIrEdHUkolagn7miD7jdyN9Q
uwGiEgtWMniPlPB9UcN8ZyH51IT/m7NIljbFCTvdiClg0zudf/3gy2cIDsFoLvP/
+Tseg1Cir2rgHbIOobJ0LKPcXkTUVueX1jh2CXLPocGju9xSyfvNVDIjZeBcBkEA
zpPryspdyyxFEuK5OPLOZ8wB95WnC9RoMCSsINr8F7GqWDImyH7REdlhDUmVAwbH
IJnpnCPGfik+QRKJ5st8zajxWTe7IxJaCQzr+fYkxJ4tcwzfogf7lnbNtcDv5CJX
/dB1mBsyL2dbqiE9W72vAgq2JPJmRuPELODedJjJVM50Li+8ACZ+x2XwWuEtd+Gl
e/SJ1gJJxerk8aPHV3tRdgZJlaeldiDBShpXNb/VQR13LXHl8xCFX+KZW+ei28i5
3mgSLnNc3hnT5GfFUczeW9kFQrtJQEq714eZfxi8Y30Le2dFKtLM4bJdUdf+/21t
uara+/bw8Cd0/JCapQWNneqIjhzsxjwnEIoRfUFcS2P5/JmMuxtm8+X6Nsvfh8M8
qsPUp+JAMPVNBoWz5p46A44R0QRvKv05gzWPRmH3mlERMBygAfqvixaSSPib+1YZ
rf3RNHyFPl5jFWO0QmQMlWHgx9Qi2Zfub0yLWIJ4QuvsTYYqNJHLAWL6ZkJk3AYA
e1GbhrtikWRvwaKXrFb1jHJFQPQFH2NsYmZfa26jAGeljZPQTVgNrg/kPrJ6PJ8z
K81lRB8+oi/hTs5scfCrtWvZjLis+YNEuyzn8bavXy2SWR+4ps9tvBV0nCU85LnZ
q6DonZ5mUmQqZwdyb2uY0QkdWwwy3Ad+5A8RQPnbwpRGuQ+JCdwwR1ehAsJdDUBQ
A5S1ESELcfIsWztSq0iP0FbJHIHToHTyVnO6stRm8pL/2F7mSjTk2+Gla766c1If
dJoQLh5xbRGgR+0H/5i/9s5OcJukVbaQMxh6sH4wYoZAIYr4Yg3iJLcjeqF9R08a
QSGRWWiDKv/djVGA9yk+lMDDPZjds65eBEi4MNL1+VEYHGxkDEOabhiyU3kj9c5U
uW70pswSe8nUOA/qkIXwVY0p5y/IxLW6i7Rn2I4wm5CF/sJ3B3I+/9whoIVYsr89
xu5CWrJV0OzelFRZiFQ9hjl48t+xei9/2CfCdwdXnmQXmqm96IKWkuWhr7OM9Zwo
NM+KHo68diO19ptppzhzSP5FqRTXdptHLXnf/mxOLBn+tJkXAGE78t56G7HKddB/
PWI8AuRmm/0YtzN74BZqyNFAoqjCp/0LjVq4YHdOIfJyZ8IMI2YgZp1i7ZOR5lhJ
/w/SphxDssTUtp3/CevqmrECU9Z5IUNZkIW/Msa1jC8ccuZ3AfG+SK9MPozU56Mc
CGVE3QR/sAaHC8SsHpGFIVQvyGX6DkuAXlJsTqTy+834MtuaiHrHDmXtsx+ySHgD
0a7krT/3+BR2ydapoTU3DBvyhqGClPopYgy0O8CjskE7S0y3LPhE7NIt1Do69FW0
KWHWz94+ZDIiRpo9BIpBr9eumGjABURt6mWRo6idEYABTGyEoff+PCLTcGVxmNdS
HrMeznXLDUZ33Qg5R1yYYXnCgnAe3q5+7WErW/dPlcGFRAfnmVtW/xNvrjDeivVi
okxn+ofjqnrTfZtYypWyHv3xtl4you+5foPNK5GSRfN+xN7r1RH4lkiU8GH+49GR
2WUciXlLZKs4/aAwRQgsIzhyWpOumMYXgihNN9ufJBheEnMvUx/fxX4KT55tyKm7
p3Id3DwazSFgrYuYyqoM81P/foh7bICa8hbP93dpKxCd/sHlF69BD3ebe6AODtDV
zHYX5OR9kc1h0fEFZgzPK0cM32bxaSqFD26LY7fxySjguw8cVju6+JCRzo909m5g
mmMI6ZSI8OXYIBdwPwiB2NGOTkT4yqNV9K7LAcvqCiV7Aj0dnJgvUELgNEaQ/b9h
LrlK77TCrwv2i+s5kX4MZpG6BeBx42zFio0uhUctoQ4y4hkF1PYYSfVufl3XPwe5
TtKA6cVNrZPjQHuLA2wjcUQRo/po3CR3/cUqy9IhHL/21FKa2e+3tcTKnulQki97
9dtWYBsJOs6/XJ0Ct3FedC3pIJS6hwSjmVi6fOdZERlYveCeLNX7TPzxOqf+jRm6
n3O3WDm80LFPuEevxtCUziRO+YCjxYzG5UDcHLH3YnSbFJVL12vWeck0ura/TsWc
lfhbezh8/GdiTqyIbOtmITLY5jBg84+Xo6YqnXAlJBhxbR3gwZM8VOVDXtYareVw
cv0FgbOtuz0/630e889boi0VnuDOgs+31k5TZCi/zyEujF/XVmmMKvn+KiQ/LAZ3
Ggj1Em4ExMjHpHizxQWewxYzxYoBlf0Iemdtwu4ESxMUQsr6+AwAywZSGKffiRZ0
RCxe99X0W3WEjQostX5brpDxG575eda6zx3d5I8sdNyph0wR2Om31CvA4tT2DOoE
GyuJf91gJTF+SJ04hoSDMLII6yEAiFVdNFTAQLz1KEyX1/VOEb5nioZL1DDylkNO
qlMWsjSOys+6TqxoxxhudewCJDbXMcTdw7YKCtcBMhf+CKpoRcK/uM79g7CfFjs1
/VoOPJJUXRmpgkafoO0PQvXtIX4U0IAyb6ekB7H5hj/B5XymX+SS2UGQ6QsdU+PS
YfWT58RrgvVHcHEDIzNGXv8vbzXJP6U1a+886PSceqL/QnvBCPAFm+HYkxnr8v6Y
f1INtML9270PtuxGmZ2aQSrYF6dNdP7VJl2LKcyceWL7w0sEsUtFcGzjFjsKtvou
CnCpPq5x4bJJLEeEpR2+d+VsD/KuUEUbgsvCJtopFX4zDDFONu51h5HqxFy31TSt
pakKb6NnFes9fI5dcNsOkmTnIdT3+1M6P8dmvGMu/zP3tcnOL29S8orOvIxmpCUE
lACM0gltxcCjXqM3Dg3iekisCVYF8qhVhRADPhRaJHepsV876S3wb7RTFRLJoEZ7
43hJunbBN1g+ej9M7qMYcWKshzORVSIn4hbm6MKMTN8Oqt8SulKQ+BDypumCa/SJ
MJ77nmBWFEGUTI7BxK0CJurEkr9zkQpn6fdhe9q9R1+j3dtoM/8qp/k8PnRqecPI
TOt0eRJBFNxomL5h+nOnkytIXf6OLyIv6c8UtC23Irhf9FHlJ0A1/XS0y9LIezje
uvDgyDWm55ypMuAJ6JnOmohLeX2j7972gGCjvxH9leB8vRvqU1nbBsqQpfosee9F
zMM56NzB+EzlFOKV4COlip7LWKwXtlR86SoDlqoatN4Cxh00aLeGowpnvAj3bHpu
QhE3wzcSSODSgKMis56rByW05Z/Z5jkSNOrnRfryzhqTVjLgB6nt7C3/q6sOldTv
TOYKeGNydJAHMoslRUN51bdmo1P5UL7UT4FK0mzWbiQtvL7A2a/J8Lhdi0RV0Azz
ih4uGBhtpKgoN1G6DRuUNLW7aK/qFlf8bnpr5vUOPoD5PzINMu69ov6LTOO5uymT
vXL/WozUvSCw4+aXjkyvCyNthldsSz1QbbmrowaNkTEtvSa9UMOMzhR+6Bc6V/YR
Ii4+kJn0Jx+AAv6KyrSJeZeMbGSmGDdaUGCveyTvnkPkNAu1gjrT54w7hw+c9B7z
2rttWlX2bWvZCvfMMgD19rQP50wXNoiBloQMxeAZd1xOILGe2m0wnQOn9OxfPpuS
a2a+HYaBTDCVZqUyfSL5VINE+uOCiedUHInxINpAYRmKa91AjzXnAVeBe4NWZu5c
Axol0uQaZyhgkKmb5ToLJVGzDHB5YhKK/6YCMIRNbDLa0/bMPZ3vdXDy8O98gLuW
W2F2B8RIqHNqGyHEc7aOX6LTYklEbTkUKmZeSur7s1jQPnx9STwkg54PF681tXmJ
2foLRjvUA7cjkRLDUkf2OYHnxHvo/HWyNI+IjQhuoYveQkALd3c6xB85TB9/v58e
NAK/C/lJAEdQFiuV3SHKZSWWv/BVQ0lyxNwcA1qLnjnwjyXLDdqt0P6oc7xKeL0N
g1swzJq3ozA/Wv5gAdiXMkcFxW2J2qbyyQhZDHt0bXnAPPb3ilRVu04v38qxY4W6
icraGnQGPQOldKzzIJi4LE2Jv1IypFhsJ3ymbq0iXPbrlKj1EfDlNOEZ3l11ansj
++joQsdRYN8YyJuR8d5zMQ65Mu9YmNAVW8NHkr4cM0QWFV/7ObglCBqNJy24XlYj
DLbFJfMPP3tINvOKEQFO5drBj4sO2h87XcHuCF1Q/XwTYEVUUYS/acv7x8zfeIj6
w0AR6oFITCG6oCs5DSx7m6LKqotGUEJmjNvyLclyGmec3fvetMz4mbhPRVq7MEUZ
We+111XeH28dvQYBecXq6618BeWB0cz+pE/5L59880hiHE4BXLqn5KZWmTjDTBJA
r0q8S2iDzie4hVq5RS+MMRXkm5nERN3gfAmHAYelLVVUxho2GTadwi+p//IWIXPW
e29bw5NU9/RNy0o0xHLfAUxYl+dKxHFb8/VZzBC8fO7J2ISB4eEayZ7j3Ph9G9Pq
Opsc1GD64xxLZPkQFJhz2mYyxJPnZJOEXMWpQ1RkplssgXK6q4xfqZCoxG/cPctS
jVVvvsT4QgEpjMmXyhXkWGAvY42msQMckCxzJ/Z1nHgF/UNf3zA2vefl6W1oS7O2
zHmXepyf5pjkcXC6KF3MFcXyci7hbAIG55w7h964eKdJL80kdh+7XSjNq1Z/veB1
ndAXdFnYJeM4xbtL3Jt3pGpNL9UhZkP2+YcMTkItiUePJzXfMwYscY/7ZIe80lPy
RiTBBWmpNkpbRl5KggU7I5XVHTLFGuAzFkaCRe5fqHw+nnDiEyTpo5FzKZLT5Ndk
5/t+cKwN+phAW5r6gA+A7fXUg4G0XeWuat45/W183Y1Ky1X6QzHbA/sLaOIcGa8H
owzFG6atDt9yJ1RZ/ms0UZ6e9PYv/8kKW3N8PINZ9RoZodxd2+LleUxlsQEQ/WBD
fMIbyKkUZQNb8OnN8XynMIa2mCTTKGV04Bb+GIoL/tRSCPZ0N2DWWCVTSSszMJmM
+6pBUiY0yJ33p1hclUvbX7lFv2H32xL2hHCfF8xniBQYZNVGCP5kdlomixPnf3sD
cuiRlDS29A7VChW9xbPUEK24s9WPdVNnyUhi0Fjo5/dE5qlEgaLPOLpM6YB2qIXt
O5wIiny2qJvrD47yq+zFS87tT6vucdtdhb5r8zMjIkLbtaNigBK5Oa+tSegIhr9+
t7RiZ9+OeSD/KWsydLis1QPqaEbS2Oj/z8niMSPrJbGQaEJ91tMtsX1ATbGNRZDJ
5moZrF1VDwcr9UqH7NNMeSlF/U2QWVTnh9nrFu06marW9kEqTzctryBkifDNOVnm
X/3xCo/soNMRLbZgGVOcYQWxktVOppHVDPpqrIHFo0/cBrdqdemBsKNGDQoVCqUE
lIHsIfmFK94tPMCYHx/GRVrgcnLZeIeeqkNQhFGMcIuAHTBBIZ0cqMJTezzlvgEl
+B2+Qw1xIq0BX/CEHapQe5zKixs8nK6WeVMyFWlvzyj3nSZwf7ZNafuXbLDkb+fW
hxmEAKl4vZbaXB0ICmwLpKIe8ZbbykHcKkBDLoEUE+8PHFmEEq7lFyHk/C2O9hUJ
ojTSwdekl8nkTYYKDpgO+q1nwBgCXvdTa1EJeCHi3zcWlPF57LP7lCZ1JapOHWlo
w8O61Dnkir0av33vnHVn4BE210ltT6ZsGh5ZItnkvQ7qhwPmwBQTF7jJABE1aHeY
nHcBo+1hf4PiuT2r+B7B+KyErYZOxPuc1324gsHTnxzLe0Rz+4ifshEzOSlqRBXs
YhI51dUREkm1K1OjPI9BVe/6Y14k9rjuwLkDllkT95aybsj+sEGyesCoqrsFmUa1
TSKpnn7KTTB0HAqlQVCnyY8HT3AXbXcPR0vcpjdXpAtO8DIsnJWcNCdRr5DWF5Y3
lvXIPY98iBKY5i4TwMp0b3ekGS7e/BclvN5YQsxSSOp/yaep6KUgvrahpMyazRh1
LUWH0Dw7xLw+91/r3JLtjn1kp2SDcrPDvmVaeT2V4EE2Xxk3TS9NE3fOwB2stnz2
9qBAGlx/juVP8yGzQ4IPOd+2uz+33/v12JxPs+N+2TrM5gMMEnj4ICROF5jio/II
srTEFHlJ4TEW01tL5krMfn86qJcdhAIvljxLVNd+PpCfvzXPsfIw0VHqDhmUSlH7
j0Am/0OJIuMfS8474p/OgLzDgxXVOXDxJmU2ColgS0rHCJJLaInSM2ZeKCTI0CCB
mhkB6NA/xpUgf5bbaO4+I2ofIf0c3xHnu7yN/+5rCKEDDNtXT2gK0Ji+x60E2n5k
E+EDBusiN9YyP8QOT1dtvUiVizSHqtLsPeTVNDASS8OcFt57fNHcIlsfJ6ypDwVe
GC+m4sHFEVnDR0nQCWAUHYNGryw7JuO4rgkVTkZQt+iTG08iHnieH2CVq3chC4Qd
zyVR0A7yve33DdamNWc8ovmmVfvhCrbNOzucMjdn03dM5NkzJLLiPpgEfLNjUeoj
Cy8ogSAgdkUHmCqUoyKh8VQ1f4oquJwM5696eXQTNLbq+Nm8JLLnjep8BCPaw/gT
ErIZvyVBj2zZ1KdTnYQOdxNVfm7jN8+dsnkynb0Nn97vwfloMgLw1+hq1AcpbCaJ
J2OG/05+znz6soq6KM6TWfWGarhpQjM6lilZsIiS4cqIJyrx6ggM5MTyM4ySUpBl
2O1bMPuF7vyyBSiFKDwMvmPpnBBd8afG4C7X4ck7Lvkc3ki5DyRmlCmzH08wx2fs
wgCi+P4rbpAqsmJbZm4tjnL6cB7Nyby/V29rKZtoXKgVkX93fr4mmWq7BksDQVuw
8lMIVHsyIo1Igy+RjO+NS4T0yCQTb/CDCeHg9yCgHcomh40zCIPiLonXZ8t41tpA
DMAFNlbPFnDK2nLrWk/5IWojIaIxWmfebOWAGdyF4VWZqmQoxv5NIwaIfegqPfXh
C/X5XunuDxyevICh2pqjY95P2Gbilv551UZaF4Lh6mvuIlElhCABLzC8lI25hNXw
tKUpoXImtn4sVDipzMxmh0ONmy4bbdRUKd9+iAdw1X+Alu6jklLaKywmeNHKU+pt
dQYw/HPTHN+MKaOpNyLD4uEejX1DLIstiwvGiFU5XRJx83UkqpYsBzg1YZ/bKmjH
KdviOAwf3OpdOihgZyR2JqQKbafwbH0pd5N2W04BAsqeAHOHdvPrHhQ7atQD+ZwC
aXXbNSTcMGGn2j3A6IOH6oeBHIecUdEEt8dLCjmiv+aueaDlptD7OoF2uY79sFnO
VNWQA3nP+WadqI4saAQtXk2sgEfiGKZ8XYuybCCNu1ocWY6ZtGb1nQlZhE/bkFM9
QHFxscpKIgR60BBPxeALWyJ7KVbdnEIBfOdApPaA6YW0XShcHBvinFNsZLCsHc+0
nY1itCcjWQLrAVV0CvmtIbD/VNB1IXyrehkXTedh37LMNAnGzKbKX6BDGeYqYa6X
nJ4yx19WGjVa/XuobAe0emeqDuxATzi2mg17KCrRZCuf8vLH3m9ZNSKH9cDPL175
vOosqw7UEKdB1DxNsboYOyaqPGIDASWeSxONvEpmbY8ez8iwvYUKnUpBTDLg2nVf
JKan3mG73BlyxANixVaffxo2B6uP/CoKRWf0NN0kweNF0CjsbwJKQJP1siHRKJF9
t74bwhsCO3I3OiWftrE0P1Ucjt3R0YOgefjBVd87xWrYqBkC62uWTRrT6JAvPpo5
8mGNSczJvbW/2z7UvYcRsSqI3s3iRtvAQcZQdzw7eumEJIx/UggmEoWMjuZsgTem
4p4Av6IQ75eMnbZvmK909KA21r/OtPot+zA/0wc+ikJC4VOBBuDMp63L6ctwcSBD
aQ2swWUl3DcBrbftMpaPhUCKfUvd65jRSDx+Qgf4wqJqYTdR4MkxJjLUtinNkW6Y
rZO+lGq3xmbg2MmV8AdmW25zn2juaZnPLS8PUshlre0VgJj8ay0i5tmFwknLcw8v
47pWWiPa5VxJKC8U9j3sz1fAy+XPqCjcHbuOXZ1ILvl8m2vjK3YuVsO/gEOfiJGO
r6csztS61QEzvMqsDxfp7zZLE1H1uprxXA5AygoVNwub9ozyKUKLdpsrsLxiwXFZ
SGzJqspGbgV1IOXmQG4MusfjtmoBD3LBDcx4b9w0VVpZbkUlZtbY/kDXEoJ0EfDI
mQgCXdYhAh/j8S9ulu2gpH+opr09+1uhRdVF2/YQ0SpRtUJ5k23sEc73PHK9KlBC
5SJysc445qZiQc/z6A5L/3pRmzwaAtcfss6v1iLIkPW3GbU9xL52KHWu8LiWUSmY
gcnmG/KsGy0keaZ1JmR4Da8qsX1AlLd0gH+iZl5N40WqnutvBjrZfnO/xSUbADql
OPA7pctTC9y9wCBG5eUpbsqVmyl/mNjx/Bu9Rer6BBbx4+l14Mef2/FZOxhASrR6
103bziy15pa2lGt0GlKz9WaPY5zBMEv0tzfXEpQRtXaaU6+7+8+BHGd7L0Htczuv
rhRXmsicWl+iNEp+Z4btUlchwPIKNFPK7FZHIu9qOyo8aR3C1+92OCAhYwGRdrjA
Trsg0miFj9dOv4fksrVsL+w3/URjeiuoB6td/Vl7/bQI4X3D4gdy7DszxUlEoF9P
my0A5TK8NY4cgjYCrunGJRmB7K2xhek2RSizjmU40EK2cX89VQNole/lgasbQsCo
SUZQ7kJerQ1jMoYUdFnSB4LkQsxDKI8908b1X1scydcGInx77KmWfvra2w5ALU7I
OACvfRC4SGdeE18OHFJKiI1Qkrerf06d2lmY0E6uiq9GBIdCR9C2N6HeJw4EqYKz
98RL2oqWaR/ONjEgL0P+uqG/80/UT76hOA0znDcuB65SLOq4UQ49YhUQDZd23dTu
UbNWHDwBEiW8YwD8dW17qmgXruq+RXw3X2yno+8gFPTF/cORY1/vZRs7R0tWZeF+
nqHr52aZno/jce2az8RO6zvaOSeh0HZKcmp2Zib4JewHj8tTU7T3bsXUEpwOsCq0
lEA1L1idlDRGuftg93uq1rLVnGAymaxmuTrEB5rO7hY5xKFOc3YDKvojHnI35OO/
BHB3ngzsxh9a2KFU2nd0H0/0Bd+2WTSDC132JHVJykuvjL8RyC18laNu/xKrLRD5
KgrEkRPaLdk9yl81WeFfozUntpp78/7sxeYMZmosp5bblF4hvABKXmCRl2rou5vx
opfVn4wHL+gFWWZs2dzG8JtHRM/CeHX+Tduyle3ouDku6dF2wgddUoDncDbP5Aif
UM5NnJH1zT+ScIAqMkZKUE8NIcjW0jMxF1WIcOSMfpzaAtBhaKczRe9rxAvJTl1x
Ytj5IwO1WKvF1p6IuFbSKjCW//yHtmEzVOGDlp+NJ+MHBDt+kweX9OdiZrA8+eMN
0q+HV1psy60ERIJP9Vj4r371DstLS/hVFxGzTWgCSMyccKCSv0/uBTP7G0TqVGM9
ckJjud5+kj1u1hgegQNFA8IwvLjHbmDThwlWEGfVBkcGit6qYVL0+sI3O0jNOK3t
5NLosq/sxZfjwU6SuESlaagAH35RAfbN/95EojIoIVJqeG1kAH6eFHpoXWhCUqc2
SKI5dMTYaWlKrDREMzpkSyZ8DbHACGBnj/PNU3ep9qXzMLFrDh0WeNBJ3T72DpwH
wB6tu2S0npfN240iplI7ykEHc6F3M0dddkU4iUWtBMF0CZNKnuuv4W/OtmBIlyDN
frmWK3Nf50eXMbus3yshSb27Owfu2wD77zcuLffgzSNGdpL1Aq4fy3p+DfjELxf2
KRfW6jo4m9/WptN3G2vXwmlnnvhEViLu5MYuv5CyW04LyevACpp9dsqEcOAZokVz
5xY0bnSESVyj8XOFh0S4EKTDqxQAC33D4LJMM5dfed62+viqAzpCy/rKX99fmFIw
lfQgkLxgPV6T0qlBXbJdojyfXxNdEyLriLg+PoAaUb5Je9onWU0q7fSEhiIjlUZv
2HFKaxYM1JFyeKO6+T1oBf5IfApnmGvP75Y1kpMYVxPPTD+KWxjQELkLvPG/Amv5
TeOJq7tT9ho83F5Rn9TBFqcOVdwGzN9fQOGAmHgBIW6KDr5QmJHoXVmkjpUV5waI
2UrObiHL3PRf2nVbT+DX+PF7VdIlNZ1W7yTxIoc2PFkOdI6ioCJOU9in15g0bMYb
SDcIJL1T4MrWegIlM6lPjM6SxczmMdO9NU0jk0eOC9lfhrcWTUlR+mrOVZfUu65/
vutv516tJUM76FwRfn3n25sjlGTT5C3NgLCl5yLw9mIRhAG/BG9xinUjI7hcNZH2
lTWBxjQaayGwojmSseFpwo48Q7IULQb+d8cFnoW0YqiiRjnCNef5xsihZYBTYq1U
PmyIWMzNpSLwWcmPVD7llSQ60e/r72TwtvkcMbkYTz162SlmJYOU9SbTbNNpw014
mL2HW2fdtwSbIxK45qxaK/md2os9+ad+eej1qFejT7iOT/Mz2/POvGtdra1/3Efu
PMnNFDYpOpXYe/rHWrJXpIlQRRKPoX1O8DKKVd0DcJTmS3Gv4LGvLXwLhNzAd0pE
oVVnV41WBalwHLD4xxZC01quQWaE33trjyqmkiH/4sQ7HNIVF+g0GBpVrsu8uk9t
Yd8YA/V7lCuiIykB1Xe9xlcv8ii6CzWBGCSKjLNUQxtsWWm+VTE5xZ0JqOtEJAUX
ODUPrfXcBkLPbCqbuAF3Eb+8UBthDMQHL5JZeypulRRxIiLUsJFsJ/9lDsVD8puR
2WqIc6eqlsNKyFw6Pa9S6JrL/x0YahMC/6g+4UgEr8bUph/RxKy0a2H+34sw84lr
ZmUtXTdvdinA7iMfY5aWDzkkl/KLJS8xbrR3imoodupkKFkqf5ff0HXflEAhAWQe
MA+bT8+gaEVfntnyMkYLJwFC7YJV178Sz8ssZKnupeOal72VnrENvs2tn4sFgs6e
esfGHrQk6rYbTTtxxdlmMJZ/aXfTr77sYZcYIif5pY0+Ng9QHJX0RcoCRR8vmX1g
8lJ3Rn6gBJkSelhpgYf2RNKZDCQ4aZSJdBMbWBZPdnn9KxCCQQSv0IqzToY2e/qo
upu4z6/I3D2AoYgpDiOuuWY9F4fcZ2HvfFtrgBEtw/uF7aAOtmMBcqdEgxoMPycj
6Atk8AsLEv6ls4mdHTHChAvtEBi5+f+R13mD/AjB0roXYJSJDmiYXCFQ6yy7l+Gw
QuXooYsvzK7qq2HQb3Bq+c+iHaCCyS1DHcne8pkmcK74TEPYizwZr5Z/5fxPYyLW
2jXJhq0jLJ58gz+F9qt99F8r6RHICeDXvOTbuiZjod+elPUCcfzPFDVckdSR9PY/
iMEOu3aePu8de6HfSHIOApVEkoUZJj5Nrd9DOa9fNDCOdFJU40ulcAUMit66cQ3Z
FjW1cRdcQgl4t1HGhTSbIeZZBC7mq4dRQV2Vhy+UjsQW9w3o4xvAYhD6WDnq8L+Y
Rxjz2l4vSc+U9DjTwRhIkrj9le206VsDfoC0EtNxEUi7oZGZGwZ7RtyBCPJxmCk6
miF8qLpzJae2VjtZzOlRqAqwGoIU7r1eWmaxP8mdcNQ=
`protect end_protected