`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 9776 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
YachDS4bpHRDzLXFQC4CtdD+ddHrS4K7VR132pOjCBP26enscjK9g7buM2ZGiNz+
2t9wy1EX+FgCtWO0OOr1FbizHJhpK628DKxboNrVuJea1KJaoEzRmJLt9mI1UcQB
IEr9b8JDNznTYvGTmVh+pa+/7+LtGxKjYicDgZwl63UkPRLKdQFA3s+NgjXwoUky
9vaUeWFA+9pAsQ5h3AY+BI/J5bh2lVoeUT/gEG61i24HSzIuL2YXt+YMU5GBpsiw
d0FbPclfuTS4y6ZNPKXtZI/9DWyiDrsKzllwYsOKMrgSxEJuc2ZA6HDNr7wibt9H
lqEUGxsePgzDLYUBYgs+G8BAlKeJMgEVYXFm/5IX+6uKHDlJApUhvYksQc8OCPuL
OjYBcPB0RLEebHeSmoyQ1Rat68d15dH4chx6Rp8w3pelJFxtP3qwvxYXYuMqmS3p
4gEs4VjpxJMRi+rZYNyBh8GxjxsQjS45B0CbbWEWT3XLHequX6MGZokvWAfVxi9U
Wk5gnWk52Yf7r2iqp2au2mrKT7WO5c3YOpIJk4eDj7fbegq56cpGjT84DT8mT5oJ
pHy8aidt+D9fBCiuQL36zI2LVJ4ZtffZGs6yeizxVhZX+tWSQn/WWQACPveF1OkE
6HKj7zBrylLRDOX/EZH0vAKjndpnNkYwTgKsv9yC0VbfhlrqmZ1raSema/DXsX3y
yIQDgTNwCAxpERG5Rq/5bYpd8cmvJIjoTXJWBQb2+zPR1RRwXT1pYgX6sz3CkWUN
XJOfGCHVgx6s7yl47LYLlQgrDQrFQNLHBxP70wLxhEL7FZcpln4DyJmKnKpPr2ii
uW1Bz/Ybxk1IhhxUXQQ+GR9nWefsjfA2lxzfHDk+5/lUpdcso/Cu6RW5PYMWWQRX
73Qpl3W7J0GfCMU6GV3cqmHOOGCTKxgJFMHSMEWUggtD6sTRVAZCaqGt0fBDAJ3o
D+62dhxdbCXgMjUoKXbqeW71b2QSrgpf3NMM84+wpozKUrmqRGDmXPwsp5xFwLvb
sp8VgbegL6QBWU6z/baDQHWhoQUhiLVwgwXj7n2kF77+EZwYIkxM1NVNegs9Dh0M
xt7gsYk8gOLnhgIN+mmYNx8TTZg3G6cFXc+Np5TJrAIYrUpYIAWe+qHjbShJp2vV
IFbNSm+I2LLjctsCn6s516iOv1FCuXaIH8/kR4IXvkfWx5DwyVfzQx0JC6CCa1Vg
MaeOKBXA++vTkF8+L96h3XpcB9p+pIeo6CkL+WBv507tJYFhxCKx5shSKs4RDO47
+MvUF8zb+fVXAOtgT5/4R5T403b/sm6bJ57E1sWFpBSnaQLJt7ZseqCguKIp0bDX
G+SBgYg6cl6+81R1GJCWfcrEnetonL1JHGvl0apOZRotCu0PN9CejTOvrqD+wfyt
2a8ztEvjWSHD0mGonz6MbcIcFuC6ol6HaoGkuoykhxzEdmiLNIFzdQYutYbUf6Zb
C8OkpFw2+gFcPUQRWGRMS+3u9YxPrfH90A6V0dKeXoZ5TOFZS6hEY9t7L1q9sh4X
qCP0nESJXr0qw3P/XGqRs7OKLbsOqmqV0qS9SNDRB9G5URGg0DkIPWQRpSPWeRck
a7sVfSnE2FAI0qWjScKStVzLd6cUGQfR6t3EjBTfnpstTtDYQWCdvQIg4yZO5YEg
ZurhAzrgNUN70RiwtSQSSu9gzzYBf46iwQpJ3FryhjnMh8iYvkwuRZTAO+hLViTX
/QU9r/9dgdq5WJruXCeRp4Xr0H7w7hJQiXTl1wI4/YVK3SKgNgMZVUqOchuzs2aa
L03cGZaODYZHeGwpx2IIHMQmIGucx03/YNYTRu+rYJI89nhzGrHJ9wJQ4jZFdedc
UvCgbuuQeknSCkKkzGTCIiDCp4fGoLCzWBMNZ9Dif2sjMyjJdUCCQodmTG67Ot65
7CJV7cZvRWEsqoXjnG0cmJsBmFu+fE5W5SFUMhwHKDXlH2eL3oFAyHOiqv4r2ICM
InGUDUi0C6NXdNyv/hj3H1/fmeiohX3l191tjZQpazKfjNPQ8nhzpvGun5Huw3LR
rNUieAPTlTS6MTsk5mg+4RO85I/BkDXwEg6l2LW50epM7l9a3P95pmqz3AEiSsFH
XLZnLUs6pGgxWOxXeGjrsbL014P+p3wDcFCf9+xEwa1ymy4A6JHGVS46X/04DE0r
jnELcDxCTinEBXoyxAkpGjEK7IUTjBUE3kmQa12/Xto7kp1U5PSQoJgmOVtQD9xn
ZWMoN3gRQq++Obvcj/WFLqSwsf19LnPUMsHKcruQRqaUKCTnNl/cMPkiiWySvG2x
jQqG+j0d2BYY6AGk7ruI4sWcsc59dOQ++3KgiRDMZrRyu3ipTW319oAsUVUMxsBz
gJCwB+pLmimCQ7WyLPq1Ii+c4Uj+DN6jOYLK3FhpwsDpAvv/SrFR1OQfN8Rb2ZFC
n3d4XuyS2OjXLE1ie2Nm0Xba700kOiIsjZgshRq0uD+GDBHmZOn2pa8re1OQotmb
6HlDGqn69bbVEHfFpn8guEDRTJ6Gb9fXdz66XfAu3njI2hSq4TUkLVrySvIPejCM
adDM2ZCqX+7Pbmsfr3UMB3rJXTpWWWDr/ARctuH0vWfwjs8cB6YmrkLF7d5TwMCs
K6SYYkUotRtgN5R5Al/6/L/lNO5pMjCpctTjYm4ZwXtqTgb2274H1ifwbUT/U4I4
Jg2+RQR/B80NfD8ly5nzSUX9cygkEVb1wgExED6A81sTLhis547hyFdcOVJkuhbe
KZgnPvOBiowzfDmj/WvrgpQt20zoC7zXyRHy27QO5Cps8a1KgXlxEsZTMV6ieNVD
hNoBzEBZ7RdUQ0NqkMoAQQhvgy3DJQu09JGYyYtK+MgZ2nzM07jS6baFQwrvPdYn
QisSMN7KhColQg45172BW+jnzXKjpdq78NXq0dJGxb86V9ZQyl/oQt+GC7saoYQ8
2/9R46N0qbqPd4udogcDP3ipY+Mx4yuYndyILzMPE16P8GdQ6nAEWv7zuJu3KGO7
i9hzJy/J5Xp24wGuasIJ767MAefrMflwhvwLJUeVLKi2+sd9BdopDQuL3CKX6N51
AJ6mb4PBj9nCqSZztijyDNLyrUKXB0f4BfEMWlzTeZPh9nCdy9U3gY0ZMnbOnV7n
thqDv75JSUkKGIJxyiyTeuL32c40FJx4fmLpO0fMGoKiZTU4ORSYNdOgJenxQmw0
E8okM9o49nrcVrmRMsbHS+VvuFA69vagobzNiLI532ADiujntd+L0x3VPBuTbb69
ADoYNNJzIgQoHCQtEjGv5xVbOFco/gyBw5hsEkXpvF/Vvizgl5ouP9Ukk1JEIBWO
hHdbddKK84Y8Z3ptSCMxo3E7VEVCDZziXVWWiaKj6+zVHoBXy3nbBqBRLz9LMSw7
HHClcwvnNHMMFZh6YdGTzeiN+WSMOAqJaxGUfGyJz3Vn0gZcaJKdFBAWeprg2Yeb
lHk8FZmb1SlSk1MKRX57QWwH9K31cfUxPYB+0ARUZt/6r8Hv+yi4PS0orkpb3+fn
OJ8ai/iXiRUj/IWmbnz6Ygr0k9AZuflEQOk/6j18CaZLsx5zJgVmizF9sR77bYbZ
gZrnuAaF6Va8GvnwXKjHzWGLQNNEtKEkYDpS4/+Mnr/Tdv8Xlx1rIrLaOg1Vsf7I
5OwyW864JbZXH5DXNtfxiE+VDlwhsky1dzpSoQP7Z9AaHQo9ZlJ2stHthspxMyIk
ls6wj7jmQpmGW26GtANX+PzQjYxVKV3eePcFHwLaFkLBy6Wsro7QNb3HZ9UHez+m
v3MoJWwaPQoNvS6VwYHsyAzsRE346AnT4VSlUaoODa+gVKgAw0HSkWBPFoSLSmvV
xrzULg/Y+WexOMIe33GD5xbfA1qSZXpxztcmMiAzur9V8hLK+5lOh5/eRI6541L3
BWfP4ndDx98hk7Rc9mdt/Uyvx8nGYO+B76Jwn0yZXQk2bWY4SuOT4XxSQ0ucLmmc
7Tcm6JrhwVwf5yPnyp2RDBu0aAdtI2/BlcypVfAytKL9w9xvE/ZcxIS7xk54G0CD
fZC0XduCHRAI5HIE2/H7JBzLjGe7KDeKV/vt2daY5FN8TuYtF+EuIc2lrrFHDQdS
B2zfTREwfYhhwGcQbhNan7c6Yv01BJjrhro/iIfcgwJH0vY9v1Gqj8RUuBHvFUqb
RJimR0KGC0RW/hLbNnKSRkKP9Erdtch9OKRylgdfMls6o1gMosY1L1JRAWQCvZFh
JSCz/LSR/Mufe1esrJ80SrA1MY76lQ55wG3EXxolKoRg+2tfzKJsHMmiY9NcWBym
fPKU6840UbkkqCOfjvUiAedAZFYNEnRx+Yt5Gp0ZIVaBw9Fjx02um9cMkx6FdKJW
q8LAu3CcsxbOyFMGHVwHSQI7giHazNfUkIwLWERlFTvFzhwsv86zlEDZgKaXyNaO
7+UWgLJorfC/B9oyQgqlN8PD5rRZd1L9KdcFHJCv41l3w5GAixBwH6I/3KcO9yQ3
pebH+upfRCPrrV8oL3/9mdkfpZradkitEZk4dkigmmgio4D5vhgybMoMQGWVJd+r
4uPlqD5zBsNUadL8WqI7OOOfQlDzRSGqNfrW2ysRQIAK51TjQHdkxf3zjg8e1IGa
KX5ll2O4kTWOqPUNLD9vo7dRscp8uJi6Nr8cnuweH/YgpQsImDaDZu3QTiE1yz+5
7M9vccT64H4u2GTF2W8/Fzn+5vy0dikITgSsVZj1ZcBcJJMXr+BwK5scI5+mVCCY
zGk92wnHH52mcy54xRa+kYksowJh04feEFqblM6DkjN/mCGjHORTQj7tU6Nnqe7S
vYzIyzMkshj0SSU8BM5jToFy0mvuXxk5a207x39jmRazKE2x4GyBLyB2TNhhaIDI
yQlpVUnuyP5BBmtC68at0AIWKbnip4qT7ogl3fagL6gXHPO7SDeha76m/4nd7ye7
ipZ92CG0HTp/g35WsSyUJVxwi8nDjoim+I8+V7JkIRl29qApE007hWDYLZZQLF25
u4zvJCAZsi7kSPDqrDPHddEEa8HTSk/tfMqbAZROvRx4m/h/E7WsLyvkBwJSnafl
MJmZJn2oZczVWAf+TSBvRg37Ls8OSorG24QZLzDJbTREv4rpGs0YnW0qj7OYsJMJ
ygh58sx/sujcVDM7Rqh3HXmQ3p5/RJ1DOR0eFxjIir/ahHByB6yql82Ww6aUvWp7
T+D2o7LWml4YepYz08JwCmZa1hKNS12RJoXlzhDCMZcp2IG7IcLPxCVfQv1KcVZ7
vKEkpwk4dZE+y7SvG/8BLKuvxNov8H7KHMESxEAv/SddGQ44V6WKYDvGM0fiqMYb
rtZdO+7ANgEyvnMfoRbRXX/9+9iXzkflRNJcRTU3238g4dwWH0EUvYWFmzTU6RUt
2fYuXby/pw4N1FS1p4c0b0b2NFPtjyxNY9ntmQo6WWwXSVo60cYmu88k2Bzx/gvc
8OyxWaCeS/BUI61416+ZbSNQz7xS07F/P2bTEwJhwM9ers2SblG0ktLNp9/llY9U
GsMmSm9lnYWYc7Z9TdGG4Ea/23U9U2ZNEjH9M61ubq9yn7SyUqHXqjmVgdm+Jy+E
tYFSWXCCmMtF279MPWmXpPPCkwSh0NuqTQtsqE95KXHknTS1O+7SrU5FuJ9j3/KT
hQ9/oxvHTtG2MWIfMRIlwDu2NVUg+qJ1bOiGGRurDCLPZ1F8g/9LiZ/D6FbVrS1f
EbVd4zI/IW4UclWfODH/1B06T4KtvUDG6xM4s458aNGfvyUkQ+aecFcXYM8G+Tut
fAqz+lfzkiKveAHi8xHnXZeUxcLk8e/0ChLOdwjNo1CVtFsAT4L+QCgBrB5eo3mR
j/U6KhPRbi5B7JlcUrX0hqLW5KyfAC8shn/1okQsixAEfAc2k+Gv9M2ZPl+4gIkG
mffqzC7F75JMvkAjHzlqs0lKwH8F/Zkh1L+sf8bE5cftWz71kT1dAXNSt9fYkqCe
JSBYktcM5OXsbXQkVCOhqLA8Ai5oPj1FSfByROlhV4ngA0BYHeb/Zxr51PJ04Lpo
9Cw+k4GnPKvnAgjIF2h3Pu+vtgSzmOjtIniJfHaRMDkhO1i4LKN3J02IRLE/2R6g
My6H9zgEeJ9NX3pQRuCwFKp12sV2fCDAUWJ8Dhm6j8Ila8lMWXXiHlf2hCm8nlJd
U2X/N/perU/axaFkPZBqJq+0az2EGuAdoAPrIDDiNGDs7qTSOGlYxMM2uDD0xT7a
MgkLfb7TeBi19LvwK73qmebnLnlBKRPebkhOCH5P1ImJ1iRrs4EghI5+y5Yye4s6
tWsOTO3ryEZRrvIFr02beeoqs7XlOWTuTfffciVLLu4rfo+q/PifBSj+mKesjpBE
bX+0TMtiV3AsiUcLHDLglmPAtqR1BqQTkILEHHzKpFbHdHNUO7lxN+gsM+E27Kh+
lDZ4ja8w3Jmdh/FEIDgjLZpgTljJAh6Dzf/R9gO00GH9/K7rNmKI/Clu/G2AJdX+
DAmoxCF6fYWkpDCJBBJl8GgnbEcyExH7GAqR83BfjoIT8bhCBTfmwRvg9IUJK/ca
s+fuYy6HlPbVEZwBFOMwHn+AOFb+yrhSEvgk/lHm+gAKcIxGuNHCXAamKvQsjCzq
RTxgOKq9YTKJJxwcdM5txpqM9Jbc+lbKBPB/MJwNhJ0jQun4fzptmEGaDCl9EMT4
oqfAdwVkbhvuTtwQIWte69K7URKu+hBO0aRV+o7Y8TJUQNCJS2tIkpQdzF42ZKZA
6ufmIRyYLYvIJI0bCzySJ+0/pTZWoW5fKxuIs226rL387bf0qJi5Pj3CnpZ0R+Sx
psMv5BfqoHQ1rxvv4KUBI0rfUUv+s5yyAWzj7635RoHH+jHN/Alcx4pbUoJNTZZ4
BlWjxd+jpPppZcqK3geh9UUTXttFUW4iadvRpHuMNO1UGuIUBJJpAcMazspNaegD
598yQD30yWvajcfrfPk2Gdg/52lpVZrNOgflSd8lRFokrlN4xk23KfFA9osHNqy8
tm/Wfm7/ZgIK7kiq4oS8gz8c7THketst68XjmebpvKMfw/9xXR7UpFH0hI1QrF7R
uOFg68HKR+sQeMCKB/BmzXEhnet10YTOgD7+a9wiec2Q97BtvjsymR2nYpG+eBMj
+jkKE7OZM5JA2SPD/S9UaFGOq0MdK1rj+szvTKMUpKdkumAUYV1Y8kXafcH9dBDI
wla/CndYaY2bgdqVyv3IrpoyzWFf+N5Zrwmk5kCGNvQ36/mq/NbLScGL7IzTcQIC
n6rwrgsRYu3hVHZ+iiO/52X/hUNFLrNc2oeDYiMbpJJwiwMnPlTohcLVifkVJ821
d9TWRki+euMrdEQThfBb6ORbS2CbMqNcQSoLSZZwZERUv1Mq2ZNlUx7hP4jxFd/1
tsVaFx5OgqaopdNIWahBcyBEMZiNxf3xaia2TS3PDVqG0PvqXF1mIy+Kzascwu0N
/ksBof0Vw0xKeSvWcBb73P3YXNJp7Erj4So+n1wtBjAayke0qAkyViCaZKj0OX0a
46N2+ZoR18Y98g+sF/EccBx0LdDYeItWiOplIoXGGCXCIRosIBXWIw1V6K3eJUYl
wmU5jeyKCuaiaWMPf1pmZrgSxip+3R0z478IaoLWNk9Ber/8IqBsyT+dWkFIonxL
IoQDX6oRskOp8SWOhtZ5iaFEAbmJH+PlF8xANTzVFecPUtJ1sMY+My4mBkJ60PGk
alSTlSE/OtL8cWOZUUj/Sagb4D+Wd2chPdNjjWV7JtnKJ4G1zcUkJwdZAVXDJ9KL
+/MkjJWP2X9pERT6BZijA9k6PfLdxAf1eHX+RyqCk2SkQkj0yeb17ORndgsUO8Vz
ehWM7luRbPOohC902ioasX+CDoPLfeIlsksmqq1L+3RcmrwA/oUznrKp34cRmRUw
1paiXfwcYBYgsUi9vG6RYBCZk2b3sNbu9Y333F7uAF9LwZ/Hw3WpUjnvh5booDRy
7ThmfGi8bwCHsfYD8NauUoATLz6LJXIhxqtwWqVn7tYth2LcB6I3o77uYLeCQKrl
3fqvFNuYj90ciN1RE6uYnPWJhghRcRE8My0RAfy/jii7c9ZW6K14fn++Sx/seVdI
dl4XrPpEtbTProvlXtK2unu3AzMo6DJDBtiAtCty+43nB4Ex+QZ7LiPwbmgcNUPy
NRyC/gqwBEvgj9yXolDJqOH7InUaVzZEA1aDfZd16Qumo+ff1FnoblcGzRflpdof
l3iB1FOvbk8oO2ezkRMAFKIaZaZ1bcgsuFXf5PQZH/BA1mE7xfYBaLQiNOsw8vsL
akMPnPKO2yPkTpr8QBVQygPr+rrx+wL+gLoLxrBjR6Flprrv8sBIAxntx+29kaC4
mWCUnnAzp6y3/EcdDC8AnjY24abFSOAubmcf2qftltx7xDAqVKp9aNXFon+aEjlg
sIC1J/CzzuAnN2dEEPqfaY5ENL3wAIZcQeAZXmEMgDS/DskrQgr7n4DIk18GGHoO
RW981vTZ86JkGRsm6MO/X+N0ZIbDgQ3ZsyCXnzkOX/6Cq8Afj9GxcONgIZ0qsCYW
ZRZlK3NL72kw/SvWNZoAC1YvXrSVkZuDlkHj2PaqjZ9X3IfVo6kbdEAzZ7mXSbYp
dSLXBO7Es9Vfr2YQeA2SolkL3efYkARQ2Puu2kuhJAmsc4Y3JzQPaSztiDdSLo5M
bCETQgQWA8ZhooY0BLwfnbgMOD7Pfq8axFRj+ceiqMv1ujoG40bROoNAhgd5vMY3
A18Z5qXj8aPAsCOKHLa+tumWTsp9pmeSG7FZN7wN1JtuJHTKDwk2egtJRjV2V2NB
mCaaniSoFy0+GRAZJiISwdXn7C7UzC7bY0SKjgmJGBfRhGo6hYeA/4vqbw8dxhML
ZTtb0TjYoKJDeJm+v1e2QwkSkVvkluHpMoaL8VY4oDWGm7eIJ1zoorfsi1r1VuHi
9Og0YfUIO+MRdxJsxzxXZwLvM+if6DULcMAmmFoLkC8iRnNSNhlVmvGdho0MFy2R
7q0wRkqgaQ2QUCr6SycVJ/tQ75GayIEMfiPzKjd0ZsHiqj4HGUaj81DwuwrR1Bef
v/xgv6mUpyZ+WwQB+tZw5K2c9XeTTC6gYkmTODEbRuG+H8OVA+ZYJ4lKciDKkGqj
Namp9scItt/GZR5I3bmlX+aMpt2oXPSqHzvUw1SU2y7gJ6VXZF1n/4i7unG7WqiO
/D4R/Z+tBUJ66eyxHVP6m26wK3Jz5fHMKMOl8Ym7T/GDvPwahhYtTEVREJNmPpeZ
nkRiNYnCKUjSPX897e8PtxVBD/oQ0zNoJuloQGiuv3oApbLCWGQ2Ko3yURZ953BS
lNyEnjXHHPcm0SUfNpRHb9ZPEFNUveaiGcEnyLp3eJX/LHNnnOVa3a14HjmNZNiC
CMUYEQ/bMyGPA3blxs/DVh7kdI5VNj7ctLtT+HDX6HXMIaSaLax/A6kqsrcKoe4u
4Z7iGEbXYllZcjElsbD3Fgenv11/jZnD4jc7NNiVaY24oJbS98pKQi69TJC7iqB7
qOqzbDuJp/tVo71jy39ggKMi9O/OOPuUL3Hc8UjLVhOF7nygGz0auBKYHjP/cnLl
o5KgzxdKe/fjTBjiVUUMzDKdtD5GCS8+Fab1G//N88OIqaQM3WQI33q2C4iSOmrl
ICyhniliFP+PcvBQ8CUTVC0hy24b+icEfG3nDxIdgFW7jpU8vnQfmowhgChcHVfB
EVAlHwFCKy3voWe/QuPHM/Mvx5K83Hh9htpTQ2eofiDw0yeasL5lDTQYDFdhf7v5
Ius/f5RqcTUYXxNNLLi+3An9WMKaL3kfWB8dj8tssbyFZNobdFmV3HEguzEvCwfx
fIyTilUsYYMkc5zUIqNcsu6T2qRbL5PeMO4DNPED7AD26WGZx/ktDL3z4qqHpyR4
KSGYAA6ns7XfjyOBVg1XlHWFoDEMrRSnl/k+zC3j4G7vfui78rXRUItGVRehEIZu
Zmd7ZNPJCG06mcgjv6CS+l2XEQnG3vnoGkj/hOWiwnw/hgOzC8m1Cg998EULhz13
EhhUfTM8V6YFsxE0AxWEgGxEIF+Rby8aA047N3gi7BedogGVFD5/HZBfazPvRiiX
o3VnoQHaDLeMCgrWhqLnemovU/37EFZ4zpCu8QO9bd2qXoo/DBaF1/ItJCr/UCIl
1VBnUGCoO4CESR9VOrrQK4s1kuZmeHF7hy0MO95+rrpEpQs28M5uqBiomQkRHarX
/c9KFq8onGM7zFeFbbIIsLhebje68AzvEnUDVnVsBsJubgflEPbyrIGXMjOAZ+IL
vp/PXRzGFi2j+/896bwHvksjRowNEGE1gCXog6KrtQwO+93QaKDJyuxfXgrAGIPd
1vIR/1YuH64+KHyJANGFjJCPivjPFB8ftN5csjhr6ZBWvBR6m8Sc3Hk5BMh3c2KO
Y4uvGZ92AdLXZ6bL+QbigbyaNBkPKGozjoIQ53l/gTMP5PhLWCnMXkt0liyWLIAl
+bnlokspY13YQhWM0jifNn0Z7dqaM42Qh/67ArKpiFcseCo3P3PVARjbezajMyPz
ujVkay1XyldLJjwiI/9UK/bsnYWGtaYTDpo0CSiVP+bDoFRtuNS4N02r70ccOpFD
RZACEYmuPkmUVR3QMwE28OjQYVm22UOfKYrtXv1rMOXiaMpZPX3UzO7MkLj1Lteg
IlWjFZc3BEsxronsFleedq3NgrMIeW4FPH3EJRYN6kus3sJvEXE+ufzSPDAbZEu8
6vB1TFmlY5GSPfUqeREpZq+fjs+TAHT+ipoKVF4pJ4p7y5nHhg9Hn9kTjCvhZwq6
GFZEy7M3oMln9tN4NAfzP6CScHj98gcQ59ZR/sx6XM6t4BJr5bKPXdkdefcaxBpo
W7Rs8gSqq6AH84sn5ZAApxRGGyuSg8kW41F7/LbtgG/x/3JG1brUe5ocWRfrEDKC
HKaMUEOP0z9NeuPkmLFE6VYBmLhBNnDnVvkJQPRZMA1/n6SKWuP5gx7KoqceTlGo
mIdvQpjMPjlufKrXcav87IrD4hW/5WYDrbTmw4xSTrT7js4f/v424HUf/fHWEJ3H
mrOp+wfFY1ORcJ/DWR9mhTT4ylvtNEBmuk8nwUBT1L3QUTQs/9ARxNhfRc9wHrEL
66xNxwMOAvK7zUm8ICZmtrjkncJFG5aamdJ204z0RGIKxoR5uRJ6H7sCsES0fMpb
s9BPHXpU9EC1PUyYbHiX1j157VhHfUsE66plt+QXIVMvVGhcX2V3XDEUs8ajR8O7
aA7Dj73pAaqnYTDA+0lak5L5t2cmTdhtAi5Nb5eZjrloPv1gWFIAtfraaqnCvWhL
3oUy/9zOdom3OXkWXkQZEEYDSs/78ZHMKvkb7wVuGp6Sx8zs8/fdyqicBtDS0xlg
m/bymWySq79m23jru57zhMFUQhBWYcnrZ7sQJ9Y9ZTT/eKYr4oTB0W8q5OJ+qyat
tGdiw60qoV3yPXs4WquA5P2o6GwdFjuyzdnOemvZNb+PCp5DNk7eSN55oS9p5GRz
5spFYH+EJ43mDYmlYo5c9sskefm5M4Ln4gn8Xa0mAWyE9xm3n4pEdeK8wEshjeSH
q3QWD36W8WEkJVH4pbMk6fp9YEjglPLUvLISs4xoH15FU7zGGkDmXWZMO/wORf1e
/9ir1fnCbFJSHx+FyOxVWhGgry340Wc/N71I7JmOkjFy4PlrDA4St/Tx3nWS6owP
cBEBPHFBCAIpPm9FLj/vk2e5+vYqzGvWPOV2vl9FJvr2HxWLanLNSwPvT3ef9f9F
s46SyjX4JuEx+fzfmscQVMEV1KpZsdPQsVvpLDDRzvQAr2P1szZQphuCUPJY2upb
C6LHZeuLUZd5NRR/+8oTRFRMo/P4kPxz/8wXDKgXPWWe4dqb/gCSAC1MdY7bgStS
Offh6YK5Op2AvHklytsvn3sPso1f1pt1C5hBXnrNeP8iZf5eQosm84K3su3nasnj
RYveIzr71EmygArBelFXozwdw5pcsFW6i0xl1X9OR83MtCEmGYguuWmMMMVV4Yl5
xXNvRcORgQs00ZoVPlImNoGCnBOhjRkEqpBo2RZxjLV1hOvqgzrsxr6Mp7cEoSOb
ftYYVBbJDYUHCS2rF4vzFoo4kg31edgi4JZeSfjAiZrcvhyauXVwirTGpXD0jZql
wS7L31W/u8ZqqGOH7AvgRC4u5fTe42RkU2jxqolwI/Z7/y3MFQmAAn+KF7mvZA1m
4GsmX7Unq44TfLy3U7P4v1IyQUPIytuH0na0woLB4AEa96ZmIF6Pd3ArGU1uNQQj
K/kWywURpaBmAfD7HuagUIcIwK3XyV9sLhLp639nIDqPSauKObnxhwbfKYgGl+dU
KeLhERW24NAHSceqLfgwwe3a23fbZnzf25PcNRvyp7PrtCN7HBqSsD93t3Vg4UpH
5tDYd4fprElPt2TlZlnCxhGroyK92mgI73Td1nVeLD6n2gjEpsrm2hcVawm2w4lC
ugasaIulfUrjxEcWv/ZlBmxLsp++lZWlSQCsUoLmCMK8wjngHCW/luaA+14YMxiN
Tj6rj6IWY6cJLDT/ffP2gjtQS+UXIbLEfjwihkq8RdmXd4y7fj3wFopDt/kbB+d0
CpZaBp2PnKZRYs24+M2GJPxTosDselp9fB80eOsgtDZc3hpmhUY2I2Pr33ZE5dxz
JK9sMyv/v7YAk18ObA8vrtb1gBPlEuSertUbmWjzoPWsMdTw1KnGPWKhpAzbwjkA
nCKIW6Rfc1s9xhDfJL0NJ9cg5Wdi2AaHXIdQGy6ANruVakkfo9HO02OcD+2Ucrbz
SNNi8+FX9a7hP0Djh7h6c8SEK/Lp/oJFnHZcljY9T0JhB6A56KONeYsuvxPErFlC
LhXisC/Y3v3PxT67Ak2WAWJnOu2yWKmtPxdkvTW+mDvhbGJ5Yd9OKBj/QaXaAjjQ
GpZsMiDHuwXSwE7KS4W69a23S0rMp2thHBu2CyfZfZQ=
`protect end_protected