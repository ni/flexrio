`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8432 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eislOGByxcl/gRn8UziAa+H
mjgbsd36EQO5Ail/O6Xu+Xx/ROMSlvuBazdeHDaf8f5b1rjPHlGu+3iGCpcm0G93
k8Sq8kYmjqgWwBdrzRzKZTfVCYH5cPa8i5k7oMJ2ddVJuLH8z38+AzMVKwzSaDtm
nKewhUtVgFiVl+Iy5ctx6eCJXST2k9p6VYLTLOLIx+gBWF7HixRrTJsJyyecGm86
+XtA68YM9Trn99Qt+/Ocs+r8CPqzhoRWPtzft/w8Y9Pb/2N+LrDkPN6LVtP/gMsn
7tpJKkAlc2kUyX+nputGP7M8fl0bNvQhp9wG7GX3WMIa3z2CRcn6KAJ2X0CK2bGu
hdxbY49W+8f5R86qEsOhES61ymANWblxKlRYUAgQfzk/6TY/CpvBEoZKu4VJ3keU
PdHKmAzSTMWnQwdzzwKbRgun2F1QV88XNqVys2bNrss8mJ+kI1jDWUaOOzz/jE+K
tZov0XwWaaxmLQWGF0FmqjBLV19Gvzk73OtfjXtWBwAtkIzRfTU793xAsGAbD7Ny
k2ksZFKoUs+kTBJRdYeLMyle+8EYk1N6VztLR3TKe/KvLMc8Ry+PSs4BEjc1rPzI
Agf6elZNZgg8gaRwBW0GkdyZuDTqu2EtkzNCyMBGuWWjFiWPBmas/b+OFahj+4qa
va+1xW32XeyGmhbA6wJqb+L2GyVREJE3QkoFc4UuyzTL016bqpAD/RjqyJE83QU+
99VuPtpld8KADETKa2LuFtJnNV3VesjNBPTfETQTrkTP2lzIfTfoKmpniHoQHVAY
+kNHul9DimW1Vh8bj+OWXLRhLGC2QsrCrPT0RwaFm0Cr3PFN5wl9hA7JT+yFFcEH
R5ZO3DQxIdsS0nPNguW5I3Ce4YwhcZzfdswu6I2JQeiDeYowsN2aps14xlquvQqt
2ebNz6lbv1jCi4qa7jZaD+yhB7zS1GFhCveLkOmIJIqd94bqmVryGkaxYzpg9bqs
nN6QC2mvY9i5aNaaIU7euBb7/X4VWHKJxVQh9S/ec1ntzR4ZtFMVIUziCwnxA5lI
sNqx0zQKCy9AoZtc5zLduogu5VedsB3PHKNRjh+56w73rVEl+SDdFOWEeQDIOa4Y
QwJfportuY4+GdIhk0rE1q9iG7V6+FNu9/2v6JI/WiXwCGWcZoyIGh4dPFOLIxtQ
twz5jk0N2ddwRBMF1q+FLESG3Vwc8HvFkO2jTaKY2TigCZP8LYH3zH2O/mjrCAuA
plMYkRGTypywEAECsMEgCl7UPOxC8fx5ux9XxZI5V9xJBzsmoLfh6xFMN7W8lrJ8
UW66r2Lsr5y3x53zog/pdXDc0FON7K1jH4tFKv9JxS6tXMnJoTuqQBBWbDxB5+7t
4IAFwVKixURpAqK2iIC4/D0weyJaVFTMlfmcCOly0oPxbidObfOhiig7pT4jbU6s
jN7YyattmJtezRaXflrS4lYuJ48oS4wjRVuL7DgieceB5gwZN1x58AgTeCIHVwDo
MBHrqvLHzoFb1oaSuC72g7qILbfeJmwlBRPTNk7sprDaHa1uY30MotiGsdaC4c2P
q43Ik0EzIUZiRa8EJx+UmKvjR289+T8Evep/QnOYoluSGDC8muH9ixeDIaXtuTYz
af7I7G1h47COBbAo347jg2E3eFDhPqz+h97tf4jJ2G/4F4mnIM2W1scdkFEb3zy+
XLVGeQuOQIh68RCFcoc0xgttSRPZDH9Six+PR+3+0p1ytxIJ7yqbEV0FwRvaC/yk
SNIkd2669zPdz1fAgRj+wnAlAogkxLfJVQLtPZJGg+V32Idwx22W6QNK6m3iCCt5
tMCaIP5j6dOOCJjk+VKeG5k+yKd3GvDLiz8MVqTeb1DVWopSlXXRJk1ACQN6z9BI
r/WXaIeb0fHFoTb80k8HZlxpDZhAtXAVSDyriKA7qYMR6lYW7nqmsKIfJzZLzO6a
aHxNWIOFLEY6laUjVHLHE8KtRmODRmHtMAKQEHj7MdO5YcvV2P5sHAClKQEswMI9
OaIWLcIviEluuDwTghH/Bbcwy6xNIC/yzFmktOnf4XbrfXxWXpJ/UlmOLulgLg/v
boRvR4z4GuJHCW3x/08X1N25+bTPia+fLgAShmn7holODljXrWArGLI30V0v+HXZ
f6KhhnJZNn3uV2ORFGiJiykahO6Z+P7HWtH10uD5G36trLSvOxes130RjJx5fwxK
MZOjaPnI5F+gUaUiMBknKM1DROGK4AANhuUhP2gXhCC1KUtv7/LqPDqkDnwm9gcF
o9tFvBt3WRHwpvG/ZKXYpchNftg8vogMyeRZMdfX76w106qyXX1FMXvy3Cucc8BK
LQzzQnjgA74AVbN8kbxB+l3g2o9IYbDrXt36NsRO1v35tpdUNMnlkC2M+VVSSWC4
WRAx9xb6206bWGLLy+Cvar6c4cF0Uw9YpDumC+TLiEYEKdca5FgQvHHzerW9lAYN
o6kBpL9hi9MxlOzSUaYPx2P8La7MuTOtRvxXVbllijiHKQN1QAYZ2uC98vyrchFx
EM+k0x9MWdH/tLN60UmppZCR3i63JXlJQLpn8YF/9I/epo+vEy6MVsZlILk2CC+n
TP+vevcg9aecAMpi+ivT/sONSthWJloP6UmFNgafg+dECArnBqTH/8fw6eUsSEGt
D/fKo/lZoJQEaW2AsDgE5MVU3jvQptIwjNFh12L9TlASaJDjALZtaa4VI9o6tdX3
Eb/zXol6g7x0A2Jm34nIPdbydWy3Ra6PNc3fd5M7uAUnQBVMOdRC4+zI/xTzTxWO
TwnvC7SKTUGncRulZ91yClKA85gLwfu/gFuyATfb9LeXzw4H+51xQNiw0XCYzwWE
jbY3B0jhdzmkK974PwUl3rQ0SMuqvJzxgxStEsnyqb9junq0+lZTOQCBDxS0OAq0
dWQaC40/rvFutkc+EgpKGtVBCdViF8c8hvovSlU0a5fAMqJtTeJoXuyoQwHm0qIA
7gFSJdv/MWPSWSJsqmUz+5bF6Ra/fPI8t56QQDejtNXvmSLzI/fCrxA7lFtBc+gR
664iTsCqLNeUgcXm8oUwvUGSfBmI5b5vnLCsN0cKcryEBlO+3U1WFeBsxZXKoaAD
bxsaEnW+977VXXUMilBXOU4B65Md+8yqTbUuxgQjoRF8qS7vF1W5k02aTvgBN3Pf
JqfjgzEeMt8/xX6QCI8vrgc0SLHeiILg4zyvpj7GgG05VLuIa768hzXdq7NoBEMY
yrcnaVagH9KKZj1JIPikTRDnNUDpflqPsg1lYYPZe3RmenVWwz4aGQs5lw4eYbsY
/sNftkMBWwRIEBk0CZlYviZleLxrogvaMqSPqFMCZ72h8oTZyLlGVgbJHWof4m71
pRam9eUFT9aeUNmdHFQ3rlGMwKt1KM7QlTzXA66Mm8zNrsK3GMujpdi2oOxb88PQ
hU0PMEKXHeRNMO3MpN7LD3/KWAFxIttpRK32GaLmT8mm9wQtTEboIuuGjLgTDA4M
EkEw7oXBrFScWCpkiTYZz6oKq6y64dV9tmYrT5kY9eTE3QnqwX74btlXlUAiqgBA
jtstKSwkPCWPS7/rl/C0s7eV30A/Uxg9L+0banRYP+FvMMQe699zYmAXHx7FBcc5
nb/uI5+bduQXC4Lz/E+UzegwT35DUfCTpBrNAcpLTyH4kEODurZNYp/axs1IIIZF
x8xQdqW3IaRk9OUTs070P5r94Ix4at24EytFtv53rSVcQuOKCBL4yiky/bae8xjR
cpBk7tZgP2qPORHBZZoYa9+26wlncuWEoiOECQ2I9ZP/WYWPvElDQxqPiZ60tyQ7
Npnx7ACWVV0HFFizgTRnQb9CIX9EJkQCYdCFHJ8dk6GNDTGVvE8HCGHuKsybNHCY
H+fdj4Y8UoUOURxm3jCwIcyNCZEe+xcorVPz0fO7m22L21lcjdEPnrXZa+rvlTMX
VpyHpR6sIAlbM+7Z9gwPJMPQwel3yMqeLnl+hlcHdNf7NTdQoLdu/NjNUJ++dg7m
yktNph8LSEc4o22UvWLcsfv4pBihuFAlImeTTGzqrnHPM15h5PP0iCuk1mS6Y9Vo
4fXmOW7Oi0grneBZm5AWyBXGuP3KyEMoABpFIwnir/PPqZObhdAKy5WhOpTcVxfK
2MOw5uZsDSeKBo/pT+nZf/RpZRlTP7sxtTGx/cgCEk/LLeCt9P2OAXw+48pmkMj/
AcmPvtXf1fICqtinOB8iVsDIVgehw4kY4z9SRWqN7xoGpcIYUMacSFTweELVo9Wz
EbElMPGwuEPZVNySD7LzBpvwbmX50zmDbFpNtWwSvm9eQ3tZi5Yz/L12Czy/3QJE
aLUOBzeLiWbHB4XkJ06ISVJ2BcUNnV/BtYOn6TEWPxrmm+gJ9zCDidbzcs3g/LdN
/ZQyaDpxoYn27nQLpbG9T9ElxM7YRCeUi5P4RNTdGeAYyJ53S+PqVaC24dvPpFlJ
dOKSf/MZS18QBDTpUAFCm+h/QBnh0ahv32aAj3LsaKRD52f4f+CAhF5PO5PMqXnE
QhQXf9tLKG938XUYRlQLbSvAQi18Z3HdJIRs6omxsGQMKYGpmcbaBk3O085tOZ4i
Ubl+M34/q7jhC6HXiBSk45rFnwb5nbGhyahdJK3zHbeaPEUKBJqa9GbeX0zl2shi
6NBF8J+suf2gPdch2Pcp69xayTGu8bofEjmK8/CeM+O1k4U8NWqXx7umCuri5msZ
L/kQCz4rARjQ4cOGuDFp8FtlcYLyPc+++rPNozo2F/XzpURc9PVff0nrHQGmL5Kx
WIqP8Saa5DWAujLNuga9Oyy/05X0jhLM/XDI/ii1noiFCmh1z/0un7kgy3JAwx+4
g87FpCb9t6nnzDSoByzuamkeVx4Pg9U7envirSpgrzJ00RRyGxpQjDx+0WWacr/s
hL5wion2ulRBSGqZ6/jdMf4/+Exqb3tXV/xqGMxhjQHIR4ahU7uqcS3efm/fd3dk
nSpXSv7wXRV9zFb2CMkRoQ5qaJXqrymShyPRfIbHxX9C6mtAhiDbC39hV+Rzqg9A
DBXIV+sn1tgDqTd9KMd/G2sUyD8HSNzlxL7YlklLq7bJQTmJbYuNASh1xo8vkOMc
6qgMM5skQQvLckZ3rXQVC0C6fHkjhnG8qGce/HChMKV8QCVjT6F6IabJO304jpK9
wkPx66A1SunrA4RLOhVXyPygQZJVRmEhPR5Q0qrI2p3iw8Z3A0i8uHbhDnRhWM9v
Yd1dIxg+J6S6StwE/ik3rVC1az9mwg/nSjNW7au8NhiYDaoAIAXIN9mX11UeYNeF
HWQkHeoJssC+GdefCwONYS2w7gUCwbzInB/WO+0Lbi2heeD5G1aRNckMVD5intZb
JqDjgKUaYBQmSa15gelhefXuwEf/1ah8s0EVeZ5DyMrpeKYpHeDLkyJY5rybfE6Q
6QVPwT6Re2FSt/+e9DUOjFgb9JFgKtp5IPsJNaHiV62iNEg2A4xPIuT8tT+WK0gj
Dqy7KbxzsRFCqJFycjNUeQVX3F0qhwQwMduQc/wDRMjCrKcyS9yUXMRuzd6jLm3E
xysgaPCtkPrfz7sJCcFG0s1yOjVFINfql1DKBBCgvyMnFcCdKimXSaHUlp3seFNe
cB8mtD5RF1ziplTUFVRoVr+rZILU69TkMvgOojtiCvuvfRSGZHSRYyEV3Llmcs/u
cC4E5eNkULq4zQ6dQNf6q5siQRhMLNzq8OyHaN0BjSfBCxvdGBrTtUEpJgZX02Vm
DqhqAlanX3PxNWIuM0xVWGYAimFHXukwXSzVl/Am2wPP1iCDxYcpkpPO1F86WXn3
osuPqVGfc9kLIxteYIVz3eOiCqj9UKx3CplI6B+Vou7csM1EFqv/5+zplrxb9y+t
UG84RZCYUg2+tgOJjB0PL5mCKOovVp6o8V+WDnkc8otenSxvYvRW6e1SZwcpzIUp
0K8DNRJmYM68lKUA/AD7AMQqYFvY1lMUwM2yc7a6CE70PCmAbdF507FC3g6Wdo2f
HfeZqR1W9+Kngi5tmpPfe0ichafyYaCpkrvJ9FBqojywq+KiQOGPzlEkXP/qEGUY
Z/fgrXANE3MmtMMVRz46ivEXat606o9JD3gBIg4DPbBL7kiWWNPbiueykCeJwXoL
CZvTc8Fbv5ebxkxQ27J/UdU5T1pUNSv+AZz3QTFDoyRhDqfQP4sHNkg40pKJAN8/
DGbvzCKmSZo9oIi38svu6+24zJL3aNRu6ZhIlHt/mKDjD5/MNW8xdqWeHn9UiUtC
jByAomudSQUWjtDVxipjHybG0XR7bJbMlsEagXZnWBW3ZrthI2cH6ed8DvofMMN6
494LxNn/7pEF7OcecNyv/p9s1qGGC2pYCjL9EVhnnpHPv+zTb4LYNRRrtsQXXQns
XCyjwrP+1jeS69A8HVUuuTF4jvZuscn1CL4K1oxeoOlASXfJc9BBnITYbj9O9Teu
x9Zf8uM6rcwLWbvKD+Qdo9Hf5tthrODxoY/KXQj/faQ9ZmddQAop9514CW7PHLhg
1abW9OuQpKkEZ+0bTJmhdySRaoiHjN1IEjLg/9w2DEG8hSCwxEpt4Q1IrbqU8s3y
zuBOkl04RcAUwqUpMHrFnHULEgiskvZ1WhJ5T7Q5PpzbxJ3zMiupkLfKl0M7F+G0
2+0MGNGvIqurID7IZQDtJfbjVIW8V/12Zx+tOIW36OtYSUBjPAIq+MXR0MbsaSBX
mYLS4lkibfrIMfjYRbbKpyAEL6+q4xIGJf9trlkgaWCTA+J2Cs+Dh9s/r4akktkI
cpjeh+OJwqn1VNOuyCdHVU+TyVGhNoittKNuX+j2SkZlHQ28BtcY85BunVP0XRw6
ZghggX+GlREg5KIidT7mnl8VnYUlamFoyy3UZEiNE/DCS9fBPhV3UzHH4XXnCI5A
ICWq5OiJ5uF8coHrUWXXj0bQ+6fUw56NXi+ST+Uv2T6gUBP0j7tTmmvfj7mydIEp
pJX+b9lB/Y6RD5y9VpnXaVMM19oOXRX1fx81jW7USFKpHQu5VIWDWyx2Tici1GOH
mSA/3Cm1p6Qus3oFhrqr3rRtlKL4BCvhj33zjON3krYbDZR4uKCId5sK+/AcK/7K
Wlpfft43lb+ezOn8q+ME39H+jOYqeqXErJuKC4/dnaiQOZjp31N1OyZC90eQXRRe
bzjKb4FOJMvuhUxBP2/Hpw0io2wBaGFPhuxUpZbtAlFbyM2Q/4p8HCT6PCVQxHiT
KRoj2uVj6lEHqullkv422FFzc2Lp//Wz+twXYPTq4VdLHM9ZEWk8fP5wP8/2b14v
eHhTzmoRXHgT5nMMdM7QfWOg9lizvA16PJYUYLstcXRgFjCl6e4AWVZDcilkBZLg
1fEa3ukJL83/p5Q/P9CdW2bOdvJGEg8jba/02/Mrxu2TksmLZWJ02tQcnbtNieM+
kyqJ5b64JOEgmJrs7VZ325OkPXaJ5Pwqcc91ioXCIINd7/wOrH4MhNiK76S7Obfp
IZxQ853TaHBGtPlvIOACDOimb/KRQNUUeFPUGAaVss59k+Z0JJIZQf+WeOFgN710
nmqgJFXvWhZ+tsHjzJBcb2TUyEXusF+El/dngNQatacoobqOO/gf9djHqxqEB4bZ
UGNE8THaoOtXCGT0toByIOZkfOmH5TdtqaAi4TnslNCAaAUCgRevmt7iP/Q4d9+C
zecGXMP6V0BAoEB4cBgVFlaUpPeuaQhu3ZvAJl+CY37Xp6wgAvvRlfdIXtYMIWOj
KT3gxDrnmBZakMKEMkVUwvKJrvvAZ7SVgeDpdSCIRcfhk239KE0mFfFqZDAHVU+O
rJc0jY/RcBzI5wL1dGuwTiwJcXqiJCXl7gl/fkhieDHF7Vg3sZxw/h9xRTRijc7T
hb1j8NnWObiZfP2fuukPRJXCVvfuHw3t6r7PUAZDhGxzc59V79pFzGMu0DTIoaGo
03T0CGhk7G7GFFYYKq0n0k7o3irJG47KCB161YVMy/HCoWP/QDj5pTWzyS7vv6fP
VQMxSRnhcEy1hicYr4jXcCOsQ951n8wxn+x3vjUJdxGczq5IXW2EEEKa06LqZ1O8
XmwL/1UbMnlEzq6mPc4rEFgW71mSOY65/Q4soQ4JLaxR+KanHXoknrkP8Sswe/aj
4KuAsvOL0ADnEbm7+SeklDnMKb3BTNH/Sfl7dbHC/JJ/loz1VsMDGtqzwfj9D2Ru
B98kBDv/SQYs7LqtuWeMkdLkim6PPvXi67EX0iErbhyMnz9Ip9LGLgdh4DzDiUhY
PQSw051gtF7Fp7nGTQ7f+BVc31N5uehfPpR5d/qzkQ1/MnxXXIyU1F3idmmyBYrw
N9VeKifqtBGQR4oXhxVBQ283vNRvOm8+bmLZqIcerur5xlJMMzRGIkKVptpSw9Q8
YP09JswPWT706kfTOQHo6s3jd01HoS3Jn1UsSgXVIiq7KTqDjoMq/bJK8to8dsHr
iLmq5V5uAn3UWmDu4hX1bDBC+M4zHzhOR1pHdBFh1yt2TsCJdm1slgac1lP25j/b
dLyzbkQrmqkS9uzs1iqsLCIumEWuCWeWe2dmjorsbDB2cdDzauPCBdEzi4WZDfeJ
Q5ydaKkWcN14T9U768MSr/w1dip+4xgM7JT2g2KYYC+xOO3P+kpOsbJ9efTmn+nI
BxbW4zTg5kkMtZ+nnSAkOtwvR0Y6ZkrBh/OgxRCa4OOjxQXF8b5uto4EM5jRoC1r
tNj8zszmrlhvWeoWXeeTPvdhLu4aWp3Ot64FrThxx/pdFAAVYQjrCg4rfVI0yd6S
ZJEmHqh31dvUkN8fJk6wlXt80UAt5bTr3W0ogWvaOgYqGfWeVCilemRl29kpAJr2
j4LhxPZ3Lf4CP2y0jm3TPPDpIZPl4oM4a7WXFeDUIqDQqs/+eudmmO2I3aVMRgHm
Gw/yooMv+svqp8+GTApfL7mWO7+kbWlBjgs2g9+KyOLHODUmBzfEZ9/9vH5qAjBb
kDYvpY2bQ9pdc8ySwkM5dYP7fCZYM7pST2yvM0Mg9wVXxk35z7rqtltX7cYl6ZuK
hMCgoMRlin/qSTUXj/SdnszViphp93wTUjEAYedirqbPhcGk0TO0PbTlhEOkZnnI
x5kqsq1x8ZpNmifVdy+W/A2WoHl62c1Ouu6lGKQxRqBL7a+51fLzUeQG/Fn14tUQ
ayep1zEC68E1e8d8OR9WXUIPCjhMRlN/WilIxcgnQoG+eAdbgLemoYXsdhK0nEag
Yp1/bNU3j8vpE9uF8eORUQl+cxfy/w1gf/uM2WGL2SDVI7kGYMBiSArLCtfTg3Iy
jyIjjdqJ27N7IQv4VB6Mf6R1nH9Qq+rrNCzFsch0ejZhDNox1DXXdOGl8MJKThNR
PaQkXE7FYjxx7Eq9P8UvAQnbPjHcH2NPDIIMZ8s9bxpdqehWasbr7NCwQ0i8bUi1
IRodOD2eX/6SKI2YXQ0v69iyvuu++Cnc7tLTFwgkT5m147vZdi1xRuBrabgQb0ZC
xhf5kkMyFsfWJC4kakmoGN6++vqKj1Ah2lnWBPF0GL32q+OcbeCyVoEypS5VKXTk
fauz5k8V6rPOpAEQ6DGWq+hrWn6wFOkqE+vjKZXdejSYfwpfPjCfFWe2H9uictEr
HbQGq/HGxtaRCnVru5DZGQibaGMe/AHIrrf5rt7oO4LvAY2TDd4xQyXLKj5APyB2
tXTRO/vBFNFfiG+FAZcLfI7n4dOFh5rgsgeuGWvaq0/buQGlNKJEJT84MpqEMIc6
vDGq04+0uzdyWTRN4VS7IDC8GCxDzCHnYiiRFMNys+8QAP78mdFGpWywNL8g6Qb/
sG3peklefVJkGqWndwLedmDPNHEHlHmBIIA9+WqeHEU04TSU7sX3ik1vc5xQaSLU
Oaa6katrcKe/vLWwBvNxKIqy071rSnOLg+jBUCJN4faYnuFX8NJlBeVJnZBmdWJ/
EjBl8F4udtzc6fUDwYF/8AdKPf0vHeJPy525vMk2xoCncbBSUSVjNy1eylGy3OSo
jQ/jV4KbSJmGftJAM313eOZTMsM9Z1PDQHrIb5AkpgHwPEwTkN8ztH/swofYcgws
6l8q10J2s7d4s6i8+quBW4iNWRK4gJMLMuX3055bMBkYNfxnqfekj9I2ZZI5J5fn
rTxklUREGPfazGADvooXgwHbA5jKoA8zicP2HeO8DEe5//S2BGQgQ/EvCn78D+Te
ln8aplKhhSP3No/Ce51sdBInr0IrVCQuu7M5Z9JKkMkMMQyYrb4v7/UQB+zGRu+U
bYvY5mzjp9ICEiyhkSwYKBNTUAe1AZSLf0Lsk2JrlmxfWp/MMSMaKUZZxZtMMKz0
sIjbWSlGwQbXUHWuit2mJ+Wbt0/2id4aglcJRT8e20QKN+XfCT61GvJ+r42MFvSN
E9ZroAQLHg2vI2qjITaIRpIHXMPAsoH5EwcvpHSVZqjyQf3x0p/Q9RmaxD1LViq0
bTqBKGgpt4RVgh8h7UI7O7xRLEtz0XkIZPjFwH4sqYvZ5mNbNNtGUwInndAfaExK
5ZDAet6sI7lqLHngPgAvNg4irWGCv1GWRZbH0AmlAwDn9GYa+paaOvQHj1WOPLPJ
8cCrXenFH//0CdccMve23kYAqRComo541gTUNUwyJ+Ai4Pzks2W1Ktz8S+rAAxTr
0PR1yVkCtp1dAZOmmuf8YeSacqQYC3baz+ViZN09ap5022ZnOqLi7NOYrpNtT774
DVAbjsWgoWSGVytKyyfT+LosOFZ6nT1rWP8NZlapdiahLSX20WYbMp0BBvOnHmVG
7TQAcdRHxM4r9zGs/byQNK3TLPdKWW6PdFW+0Oaszzxn7PEfxNJbkfC3d3QcjMDI
EpUyg4VtJqvx4zwbKjavYXiJfr+U1hlXwu6YWGaSI6IUMAAPFOXyUmJ6MDqvbULG
nx0jG8lXrE27MaVDO7AgGLWUvQREvnP/Y/TGdzOVyuYnopR4ik4sr0pTdnq8pcBe
Nux/BCmdfyO44mBPgzRpdzTFIIWPya4QLYFSpijtMaOMX82ojx4Y5J0n/ETZqmP6
8NihdMF9QZTORnDgXyG6yT9S+u2uUex7P1PLYPZrLGRKcOQEy/Hva7+lpuUyF9dT
Rm3tEvdgpKsHmUXPMbjkdGrwH7gkc67DTt4+kPQ17SKg0HKb89X5VUDyRKGIP0h0
xnx1nVISeiYkoKSAKj4axyD77ypgDc9YGtMZ2f0r1KM=
`protect end_protected