`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 12000 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
YachDS4bpHRDzLXFQC4Ctc5tISCJNegFclikZG101BG+VduvUmc14/Ji7lsAah7E
udjhBE4xkqXSTYZdF6CuLog1crgzZgmGmoWrM5FABTCeo8B7Xgp3kXmZMQJ45Fvd
C5NjPVLiRDOaS2TVbkICA4p20ZsQbqSEBYZxpzzn0+ZJNGNp4T33mvc3vGly5Fy4
dTFnBkXa6gL20YiDmtmSyF6foDqS6F3otPn7x3KWjfShnnkQNK7Hl9KYrNT/fT3J
Yv2DsQiqPDCv4+g2vHruPHUnNtNOFSVTsvoYga5LxXuHNzHbJqv8CTIFxNNu6cbA
Fwi1I/3chbsYLecWugCPdx8qtBmEDxJ7JyOuyoPKUO1kdogxijJLbF7TGZAm+C6g
JRfcFq9CQzk/UUAd6TWtZeC+PkxcRROGI7QE1GCmporetcaAmnb/gjFEoXtZCHVf
JM5Pc9P6QG8AkaFqYv6EpWtSLJ1ncK3DYX55m3p4jkS+XbAU6LfHEMyggWk2oj2N
k2H6B57Yk+DjXHGFAf7o5L1xetlf6gsRBKoqjzAEhIRQPv4dYyuwN20HsiQ2eiuR
DdtM0X7+OOfvsuTdqBDjvF7Yw9W0W/WVlqRgO8X4fo9MDPSv4wLHEhJsGNEHDE3j
yrvyVOIjAzUIw9Bml9HN89jLUQaJuKy3vibT25afoWeMMtTrzUOcfnho6rAKVD35
H4V8bULGU3TrD0cVObtpbD0BoJKXEN1S1zJnG6qC68cTIh/gtq02edAUxeFanS7I
JKFV+H+awDlyJVGP/0ZLS6vMNyq57edXB7fOXzAXSjdouj1DmcCmQcKAqQBJaoHt
s8m2eDYSLPVE9GISSIGOrqPDM4hpCcYi1RDJejmlwhYYl6R4fWFJO0Qtejqxjpi5
AbcK9zef6UC1nYvpmV+KKjuEAKmxd4s1/1yx9iAV8tn/JeyroCoLCTpEtRKoKzcc
dBwtS9MEErvy3GQPMvvz1rPWp7O4dDmdR0UbyNbqUI7B67OMqPDumsNEuzFTp7da
MCSnJwDaV5wYHoPnK4LWwlrp9E6pdRds08n5UfrXxDhya13Jt4yulsoPHKV2I0WR
EUy49t5ZBFWqz9JhshG0cQ+pO115km0py+eLjxhLqoGkXPfF0OAv2UyLhZhG77Vw
whOoG/iBkdbR2SU2Gm9gI3WPcDCHNIaKrBgQeYmpKQm/Kqpw0WhEXU9kNnp/u42Z
bMBP1W5UXavDZvWnGfuv+lhU4H/iyNUw9S/9LKtqNgJhs4od+9KUj5HGA9VPw9vT
QxCd7+aIbA05lCEcC8D1YnQuB7UhFkDt0NFJE8GtYcrKZHsr+EMoKJ+Du88doVvS
Ds5ba8bsI/TkWx78xxmgvEZl7WJfPGPfl0MJLxay8/vXcKxNrH9XRmCrtrHg998Z
ceEnG18QMQMOUSAIJfkeJPoAIjc/V74fMpGm5gWoY+7ErL+X5EQ4iz6rDIfJYwuG
OKdHPqrtcCNzJnQlkSEfHs6wm9eUsX0A+HZcmYsdZXo5iYJaDszAJZ3cffJS9qot
R7jiBDI1AgLykWHuNSmjeLf6P3s0lJYMXTljiy4IClCCfKj5hTbgDNfQZQxNuwoq
iYYKv0rjXBwU5xBC0S90l0wcVqQLuzFgMu/ojLhzNrSvb6D8CNoF4Rqlo9gt086D
PCbnitt+D6QTHZGsq+MCk/ZWND26pBJihbS1JWgGHmSwmKnld85FZzOD7q83ik/h
EOvZ9XU2DXbfpCY8RtcVBctIJsat8ntLZVh9wenv4ms1lBrPbATHiLSUygKevGeK
zvgy87rL0FdoEeXqPifng8Prqz0SvS0SONovwe5pPHABtxG8Dxw/00qlcFN3lDc5
lGVBtXtQYMMqeuN8uHBDf7XedR/XCSv+PH2P7JxxqjKXZmkmsYeUV5IhwTFAyYnt
wE593vpFn/ref0GY4WeRqIat7eiqoFsu3bnRzJzvdJU3VBqr2cBq2Kf/gepTa6k/
ihPB/NSUejYaGdzni0bB297VdWQaGO0c8Pfqp39OjyEU3zcsywm76tg/jKQ0mEP+
r3eL4SiSCoVKB8HdI6qaQ9plX8BoFN5LKgphymhkmJ3lBG/ubAyEF4Q/wyzbGrgT
GWk8YD46xL6M19Wap+y2NPjxc/gXUIVg+FBlhRmbP8fzA6E5GSj5j+crXzIym5/Z
gVwXPVYnkA/FHaCoi6pWjsnP1tNVCBrAXYhhrmbdcwwICsiW5qajK3VSUyF7EtbT
1cKlVP9pBSnK8qYJJCxuefp/SZMzx3mZ1O+Y3xN+ZQZXRucIlUaCVJjBt4qSIKPY
WOdWi3P0u8ZEdw7ioyeaHKWl8muSTZX6La8Cia12G9wlckClGMEWLfWksyE5d0HE
IVjOEW2cyMOIect1wUBQ5FnQT0cF+HJA5m+Z/kh18f31JF7VR9AVN9Ijzm1XkwXS
1R9g9WyCc7TDvzIJQ6Uffrmaa0PYMx2D10tYM0SE24DPy3oyZIJvvsqQg/GNHPlL
2AnUnvb9VcKfKmP/cEWq7t2XaM84ZKjPPemyMTwYoVqEcScH7VCNUWulUoS3iCSf
UUsQX5Spb6qQvsIdAPASkR/v+tvSwIofpz0Ch9abiRyFI/Gjc+VAOQ/WJC1k4DIq
kHs71kP/LhkjNdII1v/hh/PXDR/xKQtjppwrZEKY83zakaIFIkiMZ8zZhcYe769p
iCDDeQsAtCkAHCQOa6NPUJzo6js/tITpD/pYAtw6E8GfiLCV9POAwj0xC9ZQ9ZSP
5g4CABD3tew2WwNuShV8gCxEbniGczX2CtDoY3ogC/LriLmJRuKjxJe0FJqn9Ala
GxojFnF8ZKzhlgvmK3laicK8SM/ABECIWiwYTyV6TPB950icTvuI1ZbXjf7J9TYQ
wXTgvW28onxcvrMrtFEaJDfmn9WZk4cZwaxvO0qol9Pbyja+NaBIXU2jcCKdljhc
lJB/CNP6YwBpxnJDUyWpFBu3dVJqJCiczNMSAvka1M97WhRDBgBmoMRkOdUuI05U
rosdrpflCVrlxLODn58PDNU1BdsJzWnbkKFiNbadwBk5sfgX+dXsOR8XqTWN5DI5
ImVOk5yzButQhYcpOFFo+FIwEvxdBlCLbe9VXUV0ZP2kNQr2ZeW80nRovnG1yZ1l
I9TEnW2ZsvKPZLz1TkXVihsaKl6NKOamGn8z4D5uYgbTpIdUUWJVV2NNjaAA9ayW
HxyP6jP4AV3oxt9Wd3M9Jd5NyqCfFWk9OfyuM6FEG3mf1abJ5FSscMXpi3mm9Etl
E3LTd/3tER2gTgjXK3OVvJ0ydCxFTEHOi1YEK84894/bH9zjPvJbniecCi8dMcGn
aXoLj8CnOTH+hA666wQGVgiwoDqHJbWoEpksrKB8T+THFlDVpNlqCtKx5m1DsP94
DBjcrpeCAFEX4i/2sl8OVJzIdajzQ848CJazjvUwzPdo7wTwUOgAkInbeK+3MBCF
ZGh86NCWSW3f2eNCX0uU5C5sQRPwcwQ7vN1lrbn7cnhqAP4vt/TK5anN//J2uriW
fGcqJxwmYdILo8pDqkgmrst8rPv3NnS5COXUWX/GZSeiYSBO7UBfZDYpYTZqXCBo
L5LB6ZqIyxOm6BbHMKl5bFy1I6PeXZSWFaPbySvfec9uF5Hx7L0wQYvO+WEeq0QJ
T+QNMD7BJ+8GwZmowOySKEtQwZtUTEIciTMwAQoKaYJBUOG7uBPVqWUhOEls3tVo
TipZMoqKh9moA///DlQlZjrFh81T0DLfcDeZ0azyYDtifmAZmIpxg4OjwwyZcCK+
6m/5FtDQlUIDSEzPwZjU4tZZPsfFu+ruy1ohOJVSsXDjTKMy+EB9MzZ5Pb11SHhx
Ym1L9RnQlvLthDUdRakA1eGMVx8NFTSsRD6g9kmIJFw2K1sMb+Yydr1rXRo0QfAA
EUSlJ3fS7HEs71xzoDR0uXvhm55f7ZuZdr7BrZfmlyIxeUr8Wj7Ill5O6vcv8Pkh
Hl9eZkWMaB8eoo6Vnf7mAWElujfKq/stRX0aiz1feTbfotHJ4JThJDbCxoV8eQy7
dj0z3LT08ffJM4vgiQ88SAu2ijdRPlNyyQWa/g6JjUZ8YMbgHTn/tQuZvWuKgKZB
gmkq3UjlGn+GI1TgV6YVJ6Mu+M0vpqDaLXPAjnDU7HSRyiSXTPqYJIXNg/3LAwOY
eS00CmVoO3obn+Na5Rjs22flaLWiM87/snbXs4V13lbV8gotPpn7fzevHpSKxIz5
+W5EjZ9R6JGDv6TZ12UzM8TZGu/vLo9Gedp0AUv6OHP12r0uEoDz8OQGvm77Txy3
+vqwhB3UqyWAsac2xBDqgL+wFAtkH3RVLz2lGxVr2Hknz+wEHN7yGfjTQPwFVAJq
/kZDTIdGUb6bz/d3rJNp0U86MNon1V7Nx0KuLVy1ON0Ez19nvMpS/AatfX5kVoF0
S1nJXyfzkK9i8ERzTEF5Tc2KMgjzNjw0MyF4iODKAm9igvAoqFCHWqGy+3JUVw84
mRdrQyH1p2g33A5nnAAmNTrDQvcQ8k8XgWdMpbgHws+UYI8tntEacRkTrj4dKZ0J
PRpYgY/nimhzt61FB9HHrlPBHsfOXN8Autj0hPXKYVcjrmy8dPdcRSBuONWXfXkF
Vy7ZTDCeGfDvvUNIMFva+8+6+L6Jcb9W2LLM5Ye6OEmO6b2R5OiImMHD/TRIO1Tx
wT+yTNrhXin6Ft4A0sUbbBSvAsUm85hozeG7OGYTUk3yuF1xGclZy12yFK7vRFH6
dsbz6DjS2epAPTHuPNif7zIL4Mip8J72+mW5Dtogp4t9snbIiHITLBZa4R3SYO6E
gXxVp8bh+F5oe/Skv9c+0Z1V+SLM4hh+LmrkQ48J7DwrSoft/BQCOEVEZ0Gkx546
4YSsLvi2188vRB8f7zW+IaxeLFxsF5HziOv0leg0pp/eghWlGdYGtW7GK9iQ9qLO
0mlZRecJmpb1T/aFc98+efLEvZKKLkWPAWhf9/9yVVrOsqnli5uSeA4TABK2cmOS
xSJtAisv0hhM0UQtUDp911C/O6iHMfgYWRsxg5LV8TF9EoYY2/mII2s0jk7CR+qs
sJNx3ZVfCedwRKFwosXxJw+PZ7iPOJ+TNkDap6lgJDjNFBrrURBuJUWA6ae3TKx9
PAeYCwT9uMaFVCdZ1FXgxICHA6QZJVdbo68ep5UPfiWpt0Sr5AvmXsazAoAqnyCt
dFuXExb8IS4B/7Fr5m2J784tbjIAGFi6eDG3eK/7becUiRyarqF8dcOAeIT3YYwk
y4HoMpaXTPvQ3Ds7wOCOl29xNFROyAwQtr62jBdIbu/2rAvvOONb0KIic2dfN4VT
jR+uiNRHNc6FqsXju7vHmvyuaJoviIDP1FXdegFO3vOxW1dOHNfbws1ET02oPxfP
BpFcwv6sdFGK7SkmuObkkllfmpOW3QWnAPLEVzPzdClmZtp+/BupR38M10siRGfr
XArHei044Zj6Xhqqtq6RME+yxtHpesD7Kzu9sRB18+/HgXKloiOoT5HlLq3MjRWm
/7Q8WCYx4eAMSeiFNyTrkrTzCnSemw5KRw6C1DWMXfIk2RIgIjpAjB72IpS3oQH2
uRzPNBP9A2fPuqcTUe0JkGEj9EM8j1X1iGcoXwNUM5txXcxFy+6emo74XupAIbBe
w+DoAQ9IfiYqEhHlaT5U+BC7VsYHRmGgUsKsL+l//0YZElJPoKzL2+KD/LiZ+uSN
SNhYu9FVZYoFgIV4dYnzpWD3oWvjFGOIpS/bB+BbyYkCDc38l2OI4PYpQK7YrvW3
wNmNFt5VkvIcfpQEN2BzMKzIGFhDh+w4pqotLlXGSNqAUtTp3qNoVMDSx/JhUWff
XfJR7Pd97tjYAEdPIwRKe0qGKJBBPOzvEfvp9bsNOTq1Bn1bKq/YSUDZLnookVqS
1U4ZV0BCBQwM3mGrXaRZuOOM3Ko0Ms+wLxKVxdaM2Xc87tV3Ug4pCLKgxG3YJ+Xu
emufdJw5yimcOLd/l3GWa8DKYT9x6HLTO/57EpSxxAYfK5ArVsWaFjip2t7UrYbH
Hg9caB5Zh7Zsa9DaWC8YVmeSbbgRm0rb5k3gG0LltWX2ax1e79xRwtDTHlS9zvZs
MHH1HbKqizyqLBC0SSJXv6ano91UNz0BBEQ8VYXFvM6vDFU6J028vGYs8cU5up9w
UA/awgm31KgjNCbheShoEPBVBHsOdBWx5jz0i99CJttj6bWNN0dSADYfMQUb/3Tl
kFTnXDdHOiUT1jAdT4ZsfcqsB6UjtV8NJM3EgmWXrXSVOYtNNPTzecOr76fyhKKV
7wOitlrbc+KMJw9GWjp8GS3jHMeRuwIUpjpODx+RDZ8e20b8BmkuP5IWBfbpDLOR
2KXBeUTH9hVTqeXrjhyYB/yYifNalqy7w4iFD/QjXSPBrh6tGeOvZGyDEUi75KHi
sUReHPCQPJXiWtBqRQ6XuJaeKgXBkwPb8Pc+J7A3p1ocBYiI6xbo0ZOOf/l2jprg
k4BZwEMw68tXOlxZ6n/d/jDOkR0yl0vzhXGJLzESshGkqonKBH0tPp5HqpYfQLn4
11t7yjSH/XNpicsNNkg5D3LMXVVPPPTtw7m8izpgSTm/iM8f4pTqqAFlr8mDDBRD
USVi80ylFGRGeJJy073au1arjYXmfxFJrkdy8qHj/vbuszLAqq/YEEl+vT1TUdnA
DyS4Xspif73Y2msV4yKDhouc+mWrdbL2RqKhCDVYO0RGuSDPD6R27fEUpkxA8qne
rrfnXl8YRVoW0Mw3HhitQA9yT5gHXCqyf11GLCwfVwKw80P6M0QNLLjQjCfbvJHR
jH0wXTEWLje8yJWh1vrp0xdfTOa4y+gOY3WJQMtRG/Kx2cqyUzmKW05wcTjru5cQ
Z6rVhs3/ln8VEqD5pHXXC3laGDrcxaMn0kvGKAMhNH2ME/ICfr2aBpMOHTC4ujeJ
LZTwMmCw7s6AK1Nl/AuU/i2k5swFCMIZn5lBVsy0DTDcpVguzdlbEPWkPSqZJq/x
14HZr1TS0gUpD3tnlO/3b2QrZdlk2GxO4VhNEnbXrm1H8I3SH+EExVD7IpugSHZu
agYbECjRAqGMlr5HhUhbLRZzvFCWvNHWdKKHRYNVfm4ImIT2ZJryJGIOEEd+u4Wm
bcfMIt+AIr/J22AsVnN8l1Ucl+VCe5CQhIdoEDD4BOhpL5zXrkGgvO6sqO+efPlh
/FVpxJ5CLDGNT7+3kMTISxevzFdwJKaJ0Rb7h46OKFD4I67OsJdmehKg3JDkg8KK
Dk+93uuiwuisg9LWqxzAdfYEzKk2C3CbbceYHpzsySqPli9CfjCispDx3Hwmvc2c
ee3w9/4VR7qpvAwFV5mqWru4/4vLBQRYAN6yVEZOMkROW2GNjaGeEdowNljrHGDo
amQd0+ISDOLR5WoZzfBg5ptDlxDRyOaNQ9zWMbtMnveQhoilXz6bZUFun/bYtbYC
jAFWjLdzZriyFc/xwfPjbhVjYq+Nl1MFCEmK8LVZdjfdXl1aKae9eCa7BqXyKfNj
oFcSFosra66TsqCZxj1bmc3u/yV/gS00SvmgsmY98+uLSuPrdgWxoSRgYAURmFtG
lxei3tD/V+2vSODCb5qAb0kMyXH999LGCdqshtbG2ZUmnHzqecqKzw1+q5zRcUNg
Atoie21tOyqYYOyQT6GWlfxybrVJN7ufxL5+fAz5gcktSpZa9jc1olYNGQ/T2JLd
Ewa/bI8cU/FurWRBnc4NAJkp2fVLJmo3ukP1IA4VaAYM3b1N+oQEargoBrP40ijN
bCKN2PRiYlSBQBBqhdHcmI1gXK7zuICqnrobJP3ZsSZs+g72iIIK39vJ5TvRysqH
kjiSuwpnDtpPRUPVzmjqIORYBpLO1lvSj0ltgOjNheDFbJKhdDz6Xi3GjAIJBJjA
fNKeJKWuB3jBzWTDIL+4xwYsMko1TTS7zlK5ng5yZ9r1EHFj1xi/4rNQM91pWYxW
X4jV6WzK1bol/fj7AWoq3JzNbyRqa/u6Kl1K9n+6vivn7nxd7QGFY6y69hAikMS0
LLFPTJXyUU83sesDF7f6MrmqPG6iqOsZKyRgEXFm07cg+xeBSX7dt2I5rWXjQsyo
j0WEfUiDwIIS0NhTfRMoXoLZeI/uKbuqXQoNhFEjRDGFVfVDX+GQ/xE64bxpbkje
PRCtnGv8V2gQCW3GevP2Vur88Yl87NRJQDoE6XoJJ7PkRTv4YWLxpW8EuikLvr6D
CBdNJgN1QCUFTEoXlxRr9Z/LmVJUIvmo9XTWWxRt/BNhilXJsplct4YMKzF+XF2i
wfLhJyy5aCELeM21JqBhmtCUE30+IMj65PzAeglaS+s6QnqZHuQz9SMFDraMppSM
4Kc/k3CFTnSHqdy153SIcVt42wWcKmo00fV1KHdEcWHRiRBRyntMintClUJ+co2b
2MTI09ywz7/hWSzbUMjuTzQpI3daaIsvZuvnT8du3mpe2vQSDQT1KwGJeQhWQkn/
d9xSpyx2JL/9Ri8ZtOm1P2wAMzPE225kRoe5h4VZpvsj/dgbbsPSZQSCm/vEiu4U
qbvcMcPYLpKTYcNA8QjgLxlI7Q8sahDLm2SW+Nt+aYsACOT8kVS+Pprcpi6aDfDh
uP5jE+K6rhrbrDtd48gq7HGqh27dCZutedQZbo2MuTNFP07Y4ToLTMdFxCbypKq+
v46R9O2dmUvXzKbFXJ6l0wZvLfIkm2EQArTxig9Mb4omzGBBjALXVjKs5XBkg9zb
nDQQjTrWQ/97tCZpx6s+0kNlurfL9Vn/OE5JrarVVdOhmD2gCl7C3sPrH/MmBy12
sv+C41/t8RUx2PuH2V8XmlT6Zb+0anzBtSjjg7Rcc0YPirqOSAbRNGnF81k4BMEs
n9IZXEusz1whUZm2RabWkgKWctZmKMmQhl9ZJjLkT/JH/Uc7LeyVmQKk1V4Nz/Ry
IbMxtlSomQEDajS3JxdF9MB0hwEc13t6Hsh0tYXxkRwrcqeRO2SCH4uKMyypjSFD
952pgbBxkkjZjM4Ob5uiQKOkmBuvFaQKSk5vOHJNM46AbywwlK9Bh0VpzZGbiuDJ
VZvhFNRAlCboD/xxbuotTAOtn2wSRb5HplkbF+xFh32to6QS0zGEF3M8AA8m1hcC
trKoZIq7o+a1snCjTPOKCuq66d5AA/eeLkGFSxD2XdhY4t4i1lGyZfzboOMH0Dwb
EcXclVC4FBZFNIISPGuUdUvXN2wJK7o75N4iJRo/0cVnTAD6ouXBwI9KPTAyAkuV
3uRrfkyxn0t/trfplaioIX+dtRkn+b1bfgt0xG6UghSejw84kQy3OGSAumtgjwPm
Hd3xfaiubNQfUnNvxJTiYoE7BoHzYUO5JGSv3AnTiu8chxAareu4kOnDq+laMo3P
VD+EaNO9WMUL+4Q9Q18tVpz9OziGIQVVvohda1BN0oxskHEdOWE3u+UbYgwLGmYz
Aqv7OiZ0JCTcbnnED8m24te4SQhr3BKTfLsifzxQmAS84g1tCKCZQMgiOILKebLp
N5wpCN/7ZHkXM3WZ7LcrQfx5wKRjIUDrcj7OB8He+setf560BJjnLPmuOQuKYkLt
1h6PZLMk1IeV5SJ2tOmoCHzrp3ZKiAVB3LQX0ndz/yiki9kGWVT2a9PYnC/S7ejR
Aj1rxyllOnMhPaIt7JnDG1EILFBED8wQdDLT8LvDqIO27tZrRQp+2ZOx59dlEIOH
ZbiZViMQxwP4QY9TUIhxRPbblEyFQl3jOKcBI3gwhzE6E3QLFsKd5hFfGnRt4oj2
TYOM66QPt6vH27KSq5NgbyvU28opXDNQkMv2WtjbqIWYLG7uOt5TtoJiSbPR0hGC
OoNz8QY27e2rq+tcQI/bBG0NWTCfS3iEHhBZtw/QbOhL+yB7Kqx+yVMeNi6KksJS
vAMp8XRMfMQk7DBiUdETxN/JtxgSFnLu7Mh93tr6FVTffwDWNPHluy6LiTp5Tura
/AeDzF3JNpskcORvhDAFB0FbpTZpMXLCfXFKvthnNe2AVKNF/jUnDTqwhzV6W5ia
7BKiMUhXEBI7fDBp4BrgiNi4KZWvannJjClhMBEHauGOrYkN8dd0w6Dmmc9XYT4R
N2nuwFAZQcHE5tCWcB4wIKwB5zWTwqK77t6kQl8iIvjNe9g0pyNI2t0zjBYTuLW/
ugJtMi6TNFBtc9dyHSwaZilYAAXwyME9LxYgB77JAY8PfBdG675gUzVYfJh3Z7Qg
01RUWEqj7O6rOvV+XRjevTqMTuoSVgu75KPAD+q3S+v5194IPecJjmgl7L4qRZpw
+dcN9ef/nx9ZrgFhhJkR/ALQGTubwr5NDLvibmEVpEydwxMU8Pm4jLe1iaJLX2/s
9myMS2TXheqa7lL978pI/iAQMWt/RwAxGGKujgjeLa6SZh7jE36uACTlAjkee0iN
4qIlSRdDT4ryNGmQvtaG+pjGRvG1O/W9U5zo/IJhNuqeCOqNnd9Zlc1KSCUMnazE
d2/Ut7ZwJHgH943as0Nuh9MbaEpjR6VqzcljcM+v+kpmdYFSK+TNMd86Mq0AV0d3
83fUICNcw3QMhYwu3wi9UkuiKlUuFpZi5C53XTCoENltREGDwFM1adRcyc8k1JWp
Rvg1wP15uRqCR9TXdp4n31NmpBYD8ddygB+2QMc43zl3TRJY34M90s9N2Fk+xlZ5
dIcoQ9c3+GlaF3uCEdXFQVMXvLynjLO2JxAI/kPiyK+enn7w3uw/humnn8dkuZAG
DM6amAfziLuWwfFfhGdeZFtI7B+tACroip2jd++UVQiV80kTxJa1IQL7BCZIfBbZ
2bQCiqwL1M/mCuimkcfw/mLLi6co1KBWm4sLOVhA9WowMpRI6oai11Jcbyyj/5aj
ci5YKlzPrDNCitaZVoErwOXdYfQHG7sVH1whi0KuJ+Lk7M4rT9JllwguNAGe12Pp
Xkp4KqMQkziQvcFArRnxQmaciHXju57V0QjcqBg7qz7Yb4s2mG9k06guWSmJ5OKW
DYZ+gFABm2Y1lJ8/04ll0HDvz2lcsqKVTuCyKSecLR0QQMf32+Gr6VZ7xZ59Fkco
UKwe1jSxe3fSWllxskKe78bfkzaFuVck74icUE4FCaAxjQqG36Cki6gxHwxQ6cIS
vZRrTlYEKBYDHnRtFqUomr6xwc0VwwnwmntTFAo1sh7LY06F5GwcYrTNGpvqm+GS
ERiXV53oAoG9Fg6wK7LXspWFqOh5CH2+u4tWbkCAP66YvC1543JAEIiNTrrGFACl
nqSRX6LXEzxXjaSkCvAr+M91Z6/7qkyX//6Mkr8xEGTUVDVGPJ51SULFFhpYL9iq
atzmIAu4UbkqvO9OWX/u4KDgAPyxIqCkMc4urJbpEeUeN9lqeZ+xPdcHiGxEPOkA
dYPLLP3v8zMhEoIqzD+dsPQMQ6j61Lah4wMPGi+xvWrJWfB7g1yxt6g6qp/4F/Ql
v5xJPFV8zhZ4QRyt7K0wnm5t248QuUfpX10cocNHip31JlFkG3olnZRJ8i3bzh55
hkq2ivsGCupbyWuRHeuZTzX70XmLAugKpmLcRttDRHIdnGGYv6y2h8E6Y6KRy1hU
8/+XHE/2FyiRNvfDWg2Q6RfCjk38BhSwNShugKOTn7L+bMBX7/7mxNy6gBKe8x9o
DBN/oPYFpnv6+AcHvq9lKYEFyVi+Eb8Yvos6SbHIYDBij+bBbux3NF9SEf0R0IBB
w+1nIjlsqL2GzCV7DJD72UkoBi/6D76T4KZwxgrevaCj2PqPkYwx99FHlc1AMd18
OxjZDPYPLMlC6LDuuZjMkD6h1xQSgznghaWzvBMH9lYRiApNtKdlxy646TEn29LA
kGQSaDyRsdx0P0qQH/DOBER22n5Z50E6RiucyUV+MXehZ5F0B0OsEnXW1S+WrWbI
WN+Mmc62iOI4ZB8Ag5lic53cPVY0uBev46cx0WUJRrs/Cqt6KQV8YNHn3A1RXuf6
Yo4iihZ1Di3duJftiFhYMc59czFe94uio5qzUuYg8rO6ScgwgFct0+axv65dESL2
8Rz2wbeLFXpHvstxRuqvSr2rRT8HBklvKF+cbBQO+UBirSgvvyagnzvSVHaTE3He
r0DsNzekFm8JU9j/w46PxdbqnxgkiCHO1MhxKqdptNYTzlbeccVNOKkAe4oCSNrA
+cAKxL5p2DWv29d2lIPWVwI6y516n0CGgkmkYEpnXzVAKYy5Z333KaZy3XpMakmd
36w4C03YZllWfMo6+Gnxy5qt9YOVREc+wkMMh/8DJbtqhKTl5VpTz0s244n1Pi19
EBiKfLrxDKrRBT+mjY/5s1Wdb8nbpkBpVANfgVmc3P5sg6mUnqbHaLi8873iKhM3
6A5f1V3DzpUiHU9Vp2kMzDLFWUoFhas5TI2+RZ0OsyxycEPsTdfoGe8OeRV8RIWt
m4AxEi001Lo7hgsH2rW9IOrU3U7q7aYcYoUg8kjpFMrEl+RlUtmSKJQ/mj9Gfrbx
e43MctjatPQqPF37u8u3SD2dOYbh50nlUfqxsXXhjVKG5645K24KwG1l8MFkKnd1
qVTERI6QV4FEcyE9QhBAG22iLyiiUkauSlpf9G9csei0imAiESd4RH+SvaB4TyK/
U3GOT5SA5b+7dnteKOG/2btxUizc6b2tnLUvSCM7AAf50lMunj1lvAS4u5n57FR5
RxSs0rryGjD+NwLuIIKSjobi6Qv4ZCtN61Q2moxrccS7TFiUmoogHDkLw2Q7O9uK
/BuBriUPEFzqMsDK1TzAGLOKfoAJSVI2E5BxNStvs+DctU81baYx3EDHqQDweJYZ
aduCA7v7zpdPjty1/PLjAeGNdup2AmsESFWwEj+ALP+CUVnq5kTZ/NQ4bCAVXPCG
irO3blwCx0gb7QgU8OqqT8GbttpyYIE952LTVnrPs/qOfqkZ/e/sv1aMfcdLnAS/
m8qn2soSnKOzxJ9W2aMriLbiOcP1rlo7HgEcR0RwJ0Jzv11kumU2g3O0H+10teDe
qs8UvxG/LIeGCG0lfwUfI24woD/UTsy7/WP083N2PX6gpuEtqylSmFdqoMd+Thl4
frAs/qwO/vSUKTeVrtt9bBF/dvXBMl+OU0yLvH1nbT+FCOomopjdXVWx7bZLG2ga
QnIWVKIfplkehz7oohBxU1KpjwBJpjDmnb3j2bSDYrJI1Qq9Uja8Q9eEVnlou/Cj
raiWo+ZHFbbY87iKmWy+Dn6ZvmuzNECHdn4MYkACvBTUE5Sddh5jikqxLthrj41y
yioYMy6kfqXtm9Yt3/Ulamm/sVOlFZH2yStwZXzqKsik1ODtUVpTIV+DQTh5z5s4
j29dpAW+hCQWH6+3XG3iD7zmx8kIO42AggnJV6oFyu55rMFwfw+YMdWmb23E2fOF
t88d0HtPpbCuFbY4ePeRgLyl+iSzFvVzKtZPel9fyq18Irdt8Lw4UoQKJLpuUPfI
l/1Nx7FX182CKyxQg7M/+Jh2TBeWhqWoJARtpoX6XCM7zoycog0mnjOMEspO7vf8
JlVSWCNlN3EKf5jSN9baJV6aot+DEZ1iB34XV5nBRb9vOwqGGWvuAvnXZ9tYrO6N
7Hz1JnHXrpXcqPPSg1EtpUdEMExr6TEYSdeQh9s2EGQDDi+KbYTruY48snc6cB7U
4xoXV22xgu9KDjvE/mKMXBILIzgVoEqXaHUmGIEhGR1CfsJ+VIv+BEdNhlQh+rk7
gGx/WmvlQWRcUo5sZfAt4hutEK3GPRS+8ZBCE3SgEbS+qsJ+tT603pWpg7m8Vioe
IB+O6yNM3Xf+uGuctCYMxjbbPvLkSQJMkayYTy9J0csR/PZ6oXoBze7yFffUUMUR
M0U0Y7MoqeCzovetigdF+ju5lHu7G18vlQT8oKMhicscqcvrTPqMB/hvZUrW5UjU
YyO3atvdnZynZn8kZe949dur6G6+WWeYFdsZzocX1CsFk34m6iUWaPkemxzJMhlv
FtCXG9q/ThPV3NRezIKMFj2EIFoPQalF/cmdvxoJHzVFdG1Tfy4gcwOJFP0UD4AR
FwXu9aH8Aq+sHGSvb+mjPxwU83IXeZg5dibdIgowh/afGqCLgL96bx5C/+kui5uK
1ldSY8/DoMY1G1sQ/nMxstLiCg7BPJvcb4N3f+0ITGGEfW+n0+6WpxL/mfAvpv/o
kvTFIV/3DR6PEUzV66zngCNfSZ9EZrPI+QYBLtSM6XOEOGWQ1H/qV/3o++Hv13sZ
1zcxZc1kh2xECTqgG7PeeZoklusE7I/6bGk0BP20ZkKwePBk9XYVEJYkUum9Zbdn
Y25UwJy7qcDOda1AxZJWyr5LDUVe+F5VT7nfihoRFj4vCTGtIRwlQLDe8476TEtd
jh4mfZaalu3keQtN3QjqhRGHl06ZjZUvdsS6N3xsy+fHjGP1iM2t1fhlpq5vSeDf
+R8lopTIydN0+1N0jwzUzBnb6vU/k+QlQMNRQy8hMgDT70aAC9Vs1YEL85ZkE/uG
o3d9wSbinOSacZ6Pz8NZcIWFSjf+cUJwyKYrIB6ltJr/JA0C9AxgyZMxrhMAnmsq
xf9/msg9av4ED752KxyZbTbKcd04eI8A0329ii+PEXcCjD8NbqG17tVDcV1QSOSY
33t261/uiQWeff049l4pwLFf1U5DGTuaK6ri6twy/Ai9/q8HAUcUpJxKUvb1hkvq
b3u3IUpWFOZ0+le2G82t7qKcH+SPtkWlNRQjj0qBRzknczr3HzalEpWDHqYXOdLZ
lxXhcYOw3dYkbrReJJ+6TaUy0utx1x42BPO4cAKaOknis3DdLEvMdSuAUfZt/bB7
sO/iBN1oUc4gLCnAwXsA2fvvoP0BQ0+2NloQ/kShj85eN6IvWcXpg7AReQtMYFkC
BiapT1iFoQoiERqdPvrgLrRcnMZL3W+YLDG0Ent7VugZqni4p2M1/MlS1N9Gu7c7
KHYgSF2UKPNfboFSWAhgnNOAUXVtbSFjQcxEKwLr6RW2+JOMrHwodfHAolHUng82
atErCXREEduiOcMR/CdMFix/9scHBj2jklMZzAwdAV/OAwL7h3KTewBlbHVW3nPl
DLb2xCLfrzTkMUHJpq/GOmDkhA78PSEoBDuLDQ9RRnB4dPjYNdjWpMCvO07vYtol
iYSavP92PU+oVrQtpS8fVIMHxsWBK5mdzM1GPRkSIMz4iKeTHob6yJwshUHJYNPE
G+KDo6O2+HuDcwGC8FVZ0mSzFmrlQUUJe9gCEQZulojVnqD7faG0OK6VpfgGUbB1
GdS5R3eCWBLuR92sZyPhORmPoA3BXHMApFf1f3y6ThLCseGaXAkkVQU6cuzhuUBu
FCOfqy3PWQkH+uCXNF3JgkKx0vyh02xZlkFRKFfGBC2ofLjsXbarnQ6JJHYZufih
4Ru7AVH2VEYA8MSk6fKf1aSPVVaeBXZYZMVU7T0vAsNh8ogjA7cdZIIE2db/RVHa
dpCNRbiH3CQJ5rFGGzypE8cZ6Bk19P+08HvYZ2rZmRf0mRAPaH125RDmIVII8JSv
moFZV9eUVgISUKkNVXyY7XQZylUTJk/465S1VWvAWfSQvuGMHlXx+iS1yEM3sVYJ
lqK1sDP+rUJE5wgutFNIxwJNLT/qDggKp2119hdcuTDAfW1ShT1wHDinLUqskB7k
QoJtYRBV5WxN0gLT/TISyXrmdnnz5PuJJzucc5yRkQZ4rLJXd2Xh48+9kQ7AE0A0
ynudoTtzCqvYD0KCiETjqMBBUKnd7wxXDlv9RmnfckW8LFMp+wP47L9OaasDUIQW
cdR9cwpZ9AiimN3DCzwOJK7yWBkGW0Ptv8+eSCmxAykbSxlDy6d29hzArUgeUEi6
MOmDYp2x+ZzxBd0dDGhUUpZsehnTvi4i/UZqsy8qIwAZ80lCeyi7qiKkyEDEwL3g
CbxIeFpmjpKriZBKbEpfomSE9wmqqbJDo2O9fnRZIOklNkuyT6jp0A4JgHAizBPV
`protect end_protected