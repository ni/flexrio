`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 50560 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
YachDS4bpHRDzLXFQC4CtbN8lxqE6WQo935aAH5tNg/90eBCbCccCKX27sJX5UTf
aXBiSWqNHQapor7ao8txTP6OjHriT+g3XqJ62GGdfXXQE2WoyRoX/kMlI+Ysf5mY
uubdUjqLlIEKG5iC0joZeo83HMQ3tmkLKcT9fBEfcjK+VYL/lLrj3n7v8N49eezh
HVxO5rswkCn5xYbRyW7Y6gXGIwQ+C5ETkbqqcg7WcJaVcEoENOfg81mDr41bPyEd
SIAMzM+VYOVFHIz8aPN2MsxwQo8f2k0sQlw4OeI2vPIu0jdKhrpNEvGk5GUjo31n
rzFDRiaO6CdKbrdh5Zr67q4szsCQC+0UYG4GoTVbH0+LDG0NIYmKO5skCvv+wVxF
RjUPSHBqD1e2SUOeDf1laG8CHSX8m2MLYZn8gWqMrSCOv4sPrN2WPZPyNlh4/7v8
nWV+A7zMZIC42M7bR1XDhrb+K7dDoSDjBuUxURdEYD5Tpf3H7QsRcIhNB+0mzQwb
m2nBnHzNtv0E1bXub0Qz36lCn9E6u2uoO6Kr8iZiWT5BDvAhuzh6t8rGyPqb/jRh
YBjCAqZY4HcRrGKptRGX3X+6WBR7Yq5Kytk+R0jkvVoIXBruF0cTQaEOk7xmRI1P
E18mi/cfRQ7crpViqEPQt2W19ioVhAe2qNCPmNUfgHMNJR69Jlh1S9zoOO14PtRt
JneqzVOqIDCq1hS82dspOzd84DnrO4MfG5uozhV5QSSX2T5QWpIjOB4m2aTPMLdn
3uTcR4iwUd2eb0fzdQJj7M/q+g94lPzr75kyPoYRYR1JJ1ZQ7F57cC9rwKmxIZeA
FG65QybeRFQ8UUcAaqcsN/hKfFex+krkFTXh1aYWVCkDQcVm8IX6JDl2b9/Qfdtw
pWT0ylOxP2QiFKtoujGQNgZfeCwG/3UrhDy2rXGExN7tXo5Wmx/T1LTmxyIb5LYw
8JeBc2qB1xT6Ere20WKmnp+jErqBTRJL4B1R9nRqMubbfbLJYsgTNiXIZ3Jh1upq
uyKAZaKcFkcYMVMTgJwELV73+vmKe3VMuIzW3YE53pplNIK8OVF6McxRyVMSwCnH
ymZHLqxGaZCPWXiNQiT9sKw6eypWZj6XY1e5aHLfMLN9tG0WjJxTeX9hmdVlNMgb
TBVsWpA7uRnb1pmiP7iXZ543kCu+KW6MBmEOhFfO9JJ6hzbaHYY39IvgdtpxJljt
IydV4/0RoIl+yUd8Z/ZYI5/oPRvP42iRCB8OdkYK6Pm1Rc0vi+FDbyfHsliD2q3I
rkf+5O+XZb/g/Fm33WmWCeTqOt4LsoH2Amcz/F1u4Dx07VreEQ415c5o6ZIM6FRX
RT4Hfxmcte4VjoAZHdfsKZpIkyK8tzBJKEg9FXRyoFV0jSFO1/11IEZstHs/sPuW
G47AMluy0fhtWPFVFszWA3J+1s4QlzzBrf47gBA1OGAorsgddCQMJOXXlkrFwebZ
I47yagMCT5o9g/4NF8EagBzMB6r4uzSpUBIQ0FkaMqxa6NNrf74GzRVFZhkXvxRo
e1owAzpEynfp+8O+xRXxK/sWpa1F4u3aYCSaWPTLvYgZmZvSgJYq+IfWxR0VZysp
ef3UdLdsPzKLYa4sFo+ytJx7Aa7ZSAaEK5RzNVYfpeHI9TsrLCKY4XQKgrozvHb+
79z3dcuorlPOqcZj9Ic3j8qHlWkp2IjABxCT1wqMvnOIosJ6adWnwmvmRxae9Jre
ZbH97Ex3gn/IxAWJN+TAq7fqN3Eu7Zkzt71XkgcxughuLSZIqyr3Ub2WjtElKa11
S4Ue2Yx0ZwrckCxZGYq3C9yH8tjFu5UTsuG6dOhp/1/qdZcH5KvVxzZwRkgnnyFD
SRO0xt9CJnLw7FhXeObgPHXBCXB36InUkBjkDj9Fmldg7WRdL0GFUGsLf0bHJs3I
NKh+iR9xeqwTekJ70qxVFbldpDn09Qiaz1yT1/9ybvSM5iOpCHkW1WYKHLqDLS8/
Ym4XDkpSgNRb0TUug4xwAWDWpKgYICt0x2qxc3x4H8s94HDruuCIrNjah3hGm2Y+
TWpYa3+HWqF8pDO185SSZytVEoGLi2NSHDzQc6Bh0+MaYB42v4yI0aLilrNry639
bKsNBR57vz+Rk4mDbdjUAVx2pXz4G7YKyFb/B7Xa2APW4YaKU3rMUC40HWeM7gcH
NseJGb9F6OSavWbePgrAu1lbBklq0u+SpfyWCu5TGSZB2A4Dcy+yKL73AqKICQq1
nGGRYh/CZ3TwKBPv51nUz+Erf5XX1gEO+P6BEiU1PvTEdSRqLRm53ajADvH7Ze7h
DwuCX0lXjckCn+963JHHwEkE3wiyKdkZZdYmJ3hmQ6xq9NO/b2jjpRANqyeeEgI1
cNfkZgfmevg9Tmmz6z8aBk5w19yzJ3FFJ0zsQPrN1hii9fbJ7UBW0/4cYcWaWSbx
8oa4AvdkfO2HcqlQSVR7ESxh5QrtskwUZmhyQ89LHUPwvOyiblENZDNK8IZKIYnE
eXwL4qyI2Er4P8JEmnoKzop3fn5dKZQb0VSfiTBqlrnuhDnojgU4M2+yivdJhOm/
vX0/At4qc8+cwtrySBGmpjExgWTygFZPKYNlA1U4J80ofT/5Ppep/JW5sv4yWCe7
OYv7hBGp34eWj5HCn7WytbnOFhqw1+UJ7G6VsYBMt/kaWsVuE4Xd+jEG9zDGTmKr
CSooRBquwfAtq+5WxVbuzYA1sWr10dyKR7Kv0AY3AQlBnnzgCt2cqFASGL04CeMn
rmkGtCxwSHLhAG5fDmlA3dLGmaCnP3CjH5PXft3pPhPGz8nLZ/14UE5h+mwART1i
gOj/Y1ibbeoRkKBRGlKGXP+rGni1QHnkvfCXdldzRwTHn6LtvIu+pnu8rc3RizL6
FIWK+Llk4+bvF/NtJupeKuCsj2614XllU2q8S2AA6vwcr/zBjoH95hMlDENKjStK
jPW888oQiJQR5ilDRt2VkKJx851N2ubvWmIrMzitPDRxsg4s/JQBkahaOkc0APXS
czeYKrEsdEQVDbn88wWR/wu94RkWYzskB4ZBCa0xR2B6xCpsCg5w0VzOYrX1McPj
B7GMHOQNl7H+OBZ6p39bXoTrpsnSq3DmaliFtQ1cYT6PD+jF4wYkB761+HUUqUDo
ntVQmrQDV30Z2+9Wb7aTld5REEsPu0COI8EKFM5kv/TpqQbbLk9ksP6kudjlCrsH
L0ytoSSz0+4Ay3LIc8UxT4TXy8DhVTJ2U82PbWCXVemsoSNuNaQK8208SAxQsnoK
4ijyQn3D+4qhtU/5h9J1FMvblst9khD1L3NwEp2O61y/AqR+Ck/T6m21UWjipB2N
zQ9NhiC3K/42ftCeiMEMj5IAnt2e6WbflT3baYBZlqCGGsqI3HyNu1+SGZv2lEoA
ZnWDNBEncthA3zcsG439E9XA69y5bDoNl9jI18o0rFhJA4Ga6n7xVQTO9JoD8Z4f
UEv/GhgLAYWdAUo8RKKc7o0xkO1tuhk5VxXGa5k3M+eJ5yMM4Yp2kCciLfiE1wB8
6o+iTZbw6CU7s8OMZDV4JxDX+Tj7LKqp4g/RprZX+FNRWrYPEW20TQ+EjBHZkTZ4
wryCLfg4f4ZkVTnrQjHFXEi254hbwANoEl7KZum4jpp6a7H0sa5tThqo238CFGkC
zHc/LxgEFoxLBwBVkOefSamsKcyCPjwC/3vEUCaEeQHjUPF/gA0fM5CjUTp133Mx
k66RbBs9pP7lWfbBYn4pvZcNOn3ZpxJn/SF/5PHtyrflbxrYntjQ40RMXfzDHOwp
DYI3BYOU4Mm45R8sJX6DvMlELCmSugpaU8+p2YRyANL3cSfLBORVoJfEPOYR1O0b
m4kY1DKzhy8z9m9jrndOY75tb/E8UwpyC4a3Ydpg1J8aMMctDVgUCrPhHicXHrXc
VdgUUowGMnC9jWhiy8U5xKvMLJrW2hPZnUWi4aPP7W81Q7t54aeLy4GuU+agVGg4
oY8XkaWUBH3yUlLmQdCeppCkEYSUia2s3H79DM/RKRt5abYGCzot/uSS4rgjEbUF
TJf+TN47uH9bBYz+iQV7bZq8VPp71AVxpyhDsxLkpKmLl0+L0j18r62d5wAHa+iU
7Aqz6AWUwPxzPV7gWpDiLFDuS8NeJHisnXANUMaHVbbTmmTF7zMvw/wlbpbWVlJg
ZO0TV1moIx4FHYKqnRyoJs/KFQGvWDc/GkB234ELfAhlKq0jcdV1MEu0DEL7c7Hf
ZCB35X33hI92o3+/iUMbgxvSXdTCPK55VkY51KadBmyQ+rPg7ZUyCjgG+nm+okd8
/CCTozcv1sBzUfVLSo/qIKOaXF445xLNkcCQTm8iRs7HzswTW2uDY0Gl2w9TEJYw
S0l1NKinJUKapoKohJOhYXnemeTAPCfhDqJjuNpmMW8jaoV4h+Lsvy+fxfELZPAl
VX8z0vYEZsEyT9VmOCzL7R+0E8GM8qWfNtpjHbk+x1EpjRWvXAnvf4ZQq2skTX8O
opI/JhcHIDA5zGD4BItgHA9zzsgvHqh/z7W5tUSlXas/uEwozOzUOK3pePzqOYDH
mMF8GoVg8BIC1x0qJu2RdHjQuvFvG70V+kUyLN3e/K1+HazkIGVp++lSMblWUsbY
NpitAtVHIBnaHgiQGXF6ND3IJv5I4LcF3ZZwz5UGlewJMq5S3m6k776Z/dDA9zxq
TUZPR72m9uLThGG2qd7DBanNFz9te9ZWSU18gjVG3CpNubmZIexmT3YIr4vkAQdh
CzY83ADeukuKbto/ZzeuUBqul+117BFOiZE3hOwm+UUHIQzxFE3GHS8TbiN7n9iM
u+u8TVKXgL6Jtkv25fT/g5yrLINyIpVzfROdlXFVwshAHu2P9krq/Qen+44bl0mh
0XNo7Kso/AA/MKG0r+kuZwOKmDQ0axQToJ9Sn21H4GfIyUE77y9MHJV+c6ZL4WRq
+mU/C0qsSht1R1p+7/XlP4w/tHOOEuiLDAb6MsQA6yGJtlXJQDNQ9aYsy3X4QzCH
aP1WCgcAS2qm+jI9y13MMd19m9FzPqZd5+JqpG9T7kDMXSg604ioAgxTytXSWuqc
JPqnsQg1bq9WIiffk2mqXDLvlSbGM2Q/iViYKWZFuZ/n4aEEMdSTKtfg3PBUvYbR
3leOY9sxeFbfzmLOl82R9vJHIXRxsN16hcbaV27MBIi9s2ip5ywcF4eS1yCyU3LD
+6/2+qOQ33FaA5/j5apeEnedCS3OL2kzsGo6QCiarEv70WKB+OsRa1v3tqexEQEc
E27JUssCeGyAgLjAUZq1nYBZ3Uc94lJevjjqiAcBpvyJYES01cKhBd6xoDT27NO5
OiVFIqDVjm9Nz8TAlRHZ3orHvL/yxvHWX+QdEaPvXo0TcKM14hZgNT90VLF6tr4I
h+Q8kQsMG/mqnQ+6MX9qXHlLA9aVy/rQ1RIsk8pXjPNaZO/hVX4igejH/JOGbt5y
tccWIFkoYqjjjJbc3qmbXdX6N4n63DC/ksb2DmBvZ1igcfZNpIQTrhceLWbX8TPk
NVbL23CQjxo7feDKVZauXNUQipfShs30GHcip56BCL2TYi2VKYB2KlB0g8lsBRUq
FNuQvKzJXgl8wj2paXDF5LpkVKcCg2MVLMzbcQiJ5iXMFgmV6VaoJQr1hF/NDh/L
BXqCb/p8gJ4FVdfNdTndYJOwPNhEAJkZLPpaRgPR+De2Mf8wzTJmLoar/meo0xcf
KLS1XMCKG66oF6I+k1GlawlWtE8WX7n1YDOUG1b96dNqO2xBmR7FoNxS7r+zcfDY
bJbgYis+Ytayfm8VV6r+EumaIKfLedA2wCCUFu0jSDHQbaiRJvwbgyK8rKjekNPt
qtM5a2IKqxDbRf2aL1VHghKV5QC3LjSAq5q8ZVBzCoEu4/bRpWynop9YN3Fvs0zR
gbLfG2X/QsfWtVqYO4+elJL2cEyTF6qcNGb45g0cSgGUwvuiF/FrX7Ysp+ILU6yF
NDnvQ0Z5SqEE9r7acaalqv2jCG1kaS6s4CdS0r0f6TK1dppYQYOa2/sb95nx5Mi/
43TyERnVMaHKhu0fxuW2TsYZ4pOxIah1loi3V7v1E0P7cezOcEEH1+wopKBNjGBN
rNU776TmqpxYFodRxvRsoyEvzShEjxU7A1uDHyjVxX1oWnjdeoGIXSSI9tXnvZxq
NDv3T1qyDvGSSSt1fSVGGPWp0ygcYgZhDWa/mukkPE8aGTBlxUIAQNi/3xpzH6IH
pAwECq+h5APPlcPFVKwysqvgHjpNcDuXfJvfE0e3BEiKyy2Zpgi4SHQkzI1qzuYe
NLg6csOH5hnbunk0qUceLcYo2S860z3LXNKKud+Sbfgca8lvIlyPRolafyA9fbBK
4QxnjsmK9rXD08A5H2BqagFbuT/nekEoFJrOw4aQSoYr0VamRfdsn1CMB6xXDv5W
7uMhtf7KOjvDW6AXRUSHhDi7Qs+Jj8RWYifTmi4LjQcNYhPZwb2dwuPSDtSXTgrp
RJxA0jwVQ0R3Oo1tq3hIKYZ+7CYCPtIl+2PFFXLzdGGuruYpeTyAXCgYiacHphk8
IZvHZCWtY0VPUZDEKnXlU7nsgQUbR3pr7rOpUEi7HzqkwghiPlwMrwKK1shI3agj
pVXoFgAJWUkvAq5caAuqJvOhh4ArWiFUKfhSs911LZrjdVxYwgNNiqZnAh2XXVBh
kF4w+7RbrvzwHMDFHvE9O/t3eI+JBuMCHtqhOIO34rLEg/0OavkJcpHrlTJTmi5b
qhBmY0UpKOPgxNjz6V64XnjBJGFKWRSjIkNHHcFGb351cbGUIRM6otwMQPbY5NuM
47KO5MdlT7IOm2bFEMxxJqCK6BWG5XLzA5frMTwY/F+vA32igdMmiQsPW4JoN69E
s8Qln8MqONi/i0eRmPgsYqSgN2845hGcqTO0SHvdX30VglnYKs/jupskfRH5SvzU
atX8rsUcjsFqSJc0qonDi1mGdEgst6K9kwZ3Ixolj4zPV/KPwKCAdmIL5tl+uNt5
bNmkXh2UbbdNF4bh/Y6RuDc1bjnKUx692qcH8vYRb3Fb+oTW8MV11t7YykaWzZ8D
N8YhfIkgwaMMC4Cllk2HJcOom4FcNCSAKSYWiMhVx0w1oCNg1FsSjOYL8trmqTBc
MJBXTdkNdgzjgpI7muRvrYqOOfYsjJm9G097jCBMDHymPWsNDHPq1e+5qAfp5Rjl
3TW27TYNaD1c8l5zR7ilft1DJfSx+bWmQlsat1iNISuqXXFEiJi3kC/NVPG8F8Ct
5jezNspxbyKvAiKY3Q+/OjLmcznsqUJu5N4e43Mo2hmptaE3a9Im8P6b4+rJ/t4b
dDGlRZSzT7m5LxGYYpTShPigD7QuqW5z045OAqTdLFO1Zs63NS1X0EPR9wUh6Xsq
CDWOy2vNk2BSS6ZRy2lLeWaKgx+D6U0ok7z92+IA77T3Ac+xzLWncyVQRWxIf0c0
eH8Y/NPrc9lM5BZjX4Q9x+IBj0qpCKiVQPWsmS4kNV9cSB78M89EqwQd9pz99xXP
jkRMhqotuzc0w/VIabkMUiShuGcq+wzG2R9Jvzs+35gp5tFtFI8rfbmPemquV8bt
5WU2sZ7VHsyJwZKleBT2hTaZiu2E4az//G1XbgFd1afHIGnKzHzsYPF50AOYnPte
CRTn9pEWDLs+vgp4WKV3/Kizd1s0JoPnvdXtEPzmuxxsAmq9nslhzscXKth1YLmF
1D0bsXycwDfGtpbh0AZ5J/pnjITq2dBtVSgfRJSlyu5coo0RDIj9MzghLQwHpdr1
tlpwA4vgj4Aynal5b5sDiGRqZEl639Zk6I+i6J8zmRgNhECOxE/MucYApaRikvmu
gsmyK6sHbcHQH3JrLhrRxOSImeCSEZnxMi7zElHtADZ0bveX+lpKAmgMX0f9ryTY
BkvU/wjeftQG3Tlgnl9RYaG517paxR6/Shsn9xroiquJcID2CultbckxErEQ8B1K
eYNzutQA7FrhUuPimexwuHFtbo+IO09ULX6YrwB7ohpw0UCAKT/iw9nLj5WhhElW
MqfXbUdSPC2POls9gNuMpTV/Qp6oNA4oEsG1qQsJ0ssZ8yNdI2qqV/cht57HPnxA
+6v5arlMBqQTWMOzdXKEWqjZyw3IStEj45nkcmeDlHukaGJjdQR/PEC9749zaIkT
TEqDR8QKS/XoosQsQ/V06ChS1WMFQgm0HgeoSXNZYup0PnFgc7M3wI1ROlNYr3sJ
3SFiyShZiuMaagtB8YcvljVG6mkD4WD62nkY4xWYBTi31cq14ZrdXTYI8LPBWAH9
bnviWgoa6lJyRGPkFvduPt/E46frGnGrT7Qel7ilj3PsONrQL37RJ6L/SXBLN4I+
Xwzg7ZJS8rjVshkrikO7QG2nfvhqIunYvyk061pDQAQk1NV9buGiLCFQ++gnoWaV
eDS/1jkfpp3nG31ygTMiQk50fJ6ZArue4kRX24UXU/DkiCS8j6DUxDj3xgyVKWyR
Tt1eaqXq0JphRI7iL+dxjCvNyH1/j5ZGcZmL8Xs4hNA7QmAFpoXoanVMbevbPn5T
ZEQpUO9WGR3sOKQmPCAHjsp2j3B2I8Yw51FqAgUI1i4SOLXUpIl6QMHCP0MLnIpq
L2lI21Y2xwq9poof2PAEZehuLOk0o5faiUxwbEbfw9cS8v7+4BXrsYo+hhQO4FES
w823bcowJs9k/F2UAKjAw3WRaxfTibtr3HohYpty8gJLbZHE6ZPnj0B+cXJ+qE0j
o/XPQJhJ+0peAo4FL6Zs12KZDCncJNRJ+JkpAoIwbIsS6McwemdBopQLLwrd1DBj
kIYAlY/LLroT/waTV396ushB6nyUWGR9l52Jxk5onpwwzQOhpaXMztgIw8WrGKg4
s+vZLbDqJxbsUGQlKOR/VvZLGAuL/dc6w7e2tJ9u6eUL6hLsG4Bjv1pMyYYVsfK0
HW6P0MDUSaRysQ2ppX8545lvIjq/zMg0XNecqH//Oz2rXFP06efyCO4tCRHWRtHm
08a3RBGW8hC8Txd5RWV95zKVUO4i9DsO2Ep03vgdgf8alWw60gtrRrTPj+3pVWKQ
XU1CqO01ssebVMmI/JzlZnduEnsqf3GB4NmSizO+y1tbZ/ZnnUdCxKC35CvA5F8c
gFb9pTblKEnTHi5rjsi36/C6DXoT25O7SXwazXV0wv4XBBqwrWJYJRqG/mw2tqBj
ETSm+rmiqTROYmHfabkqrIGsBoukZ6Jd3AEOHvWhIdcKYgaTRJydwG+4cCgJYDEH
eokhs6sHTvIR/cRNGpSJLTLrxGTGo8PIdqVs+IiuhZdInDAUyN5Euy8DwvC2F8iT
6ARcNC+oAL6mNquDMxmX9mr8Dj+TTGIN+fXmmR+wHGAa3dMsVnRuxj7AbYHcZFfj
8O58PW8MrsJvkrEa5wPOcsww3nJgHSWNaS/H0Uk7/QqEIv1Af42irTZKZFijHVUo
3MTecdVJipE98dYAL7FKQIvjz5bO+xESAa4aSQbU6zvCU1m3MctR8UfH4G44bbzZ
vZQ9FzjbYNkYO7k6oHFPso1cGXjYdJkVVseXUjb4LUvZXxFPeOHUU4BV605vU+GM
SV50m7EGSF+ekJtWeP06A8gekYJWjGoRXKskrWQAjq5kMBgKG9Kjn1a0ZicxVmBD
MHFR5V7uQ3VWZv1iUw/h+vFZLJHXC1C3CEPqtMD+MYGf3TVsPoILKo/YrQYMN3W2
53n7USembcoLjWL+ml8LpRbT7Ub1o0/212T8uJyqxX3cOtqF1KHhjF7LX1WS7q2m
UYrVp/cOZ9xx0K+bceI4LE1b3UKpYkbHFZUcFL9TkY98Sj3nxxQDNN8cIQWVfVvS
7LlecchEW9lv2WxnLwD/s4o61GOd+ExWt1uMn+HZSjNosyhhhj82Qg349B1GYqDx
WiTT0/gYlOMNkzRqZuor6mNT4wDggI04IphR9dCyZu/UnwQ2A1GCIMEeqiBW60Vj
QTu8+7x0+TYOAX2+dqjr5ADH8P5PXP6yrWqLdDXYgu/eY41dGO8z1GFwwjb+qC5K
jyYgP9g55b1xsFC2AIDhRkDmjY1zOqOCoUDva/1q5slSjzUfS1CHYIH35SmtY0ea
VZhiBlZ/LRvcx7XR2KfHozgzPMfibgntMJW+M46KGniB1JzXDjUB4ECJ2waqtF5y
zOG3hKO88P6/W5NJC1QPBcYIiQ5zxv/0Ef+cZu4KFQJ//o1qSSlZz61K58r48l3B
tjI16ye4O4pnWVG58iAms/AFG+UZQ5TtPus6FsfYVBQK4udt5bsMAgwgGUJ4l9Sy
5yHDzhIgsSTBeihkxmaVU9udc9uUDzOGebfE3K6yLrk3eFo1ujavVu1P0uvv+7rF
kRjXR3XP2Yrkcpk98ITIeSnBgfg1w2QZG48vrwePZdOGHkKLIonXCKBsJL9ltR6g
EgN/3Ypt4+mwyWjbBbiU0QRk//eSkgs0yfoWHR26b4+wTTEKcfZIItGqANT5f35V
VV1ZuJN+7i+XdxgWtR8+40KfuDv18wosqS8py84Mz0vH2t2WwpAETf8211h0kcKq
iRuKB85RTyg5aoiN0Ot35rIfx2eZJWfXluwEDH/kZlNDcwcoRb/tjgjT+uazUGn3
kvcFNJWv2Z19GIauUJAEjoVVkTt1I0haGgoiscYXavPFcPBYrkUk5jOz4nPxDBqX
yrQGaU8LJMPgRebOIOhoU/ltj5RDn8pl/QgdDCPlsKrOPTGJIcKbXcOsKW6F46Fo
XdzHC3AUyksZECUNmd9w4melmXhybj4LD9WNLuuSmctKpzhMp4lkyOvpoQs2Pg/K
URleH/7hPXxhVv8jPHg5vlx4KN4CYQI9VNo8289CuDePQEjTd5FyKX+P+m/WMc+2
mtLSeYGkzn19dvDLVaGtitZvYBdh47MESlknWfiISkU11dYpK7jqvo4SyBEK/Vxc
vGY9qzwfZafOUfE7FZhq1BUQGQXDeogmIG1bZKsombxYyiIZkLOYk5ZMActqkms3
gT8axULZTtsOJL57wu/Tus1Rwqv0kFwert1hXlTIhfBz3StoEZm8pPkLVNZngD+b
rI8iE/CRt4Y5Mtd+k8+mEMS/UYrP56kUm8sD7OZVNqJwqc85xz0sJ6UmzI6lxXZm
hs3jvp4TX3SxX/YRl29c/k6ESXP1LjHvN0EpiA13H2sPzRCIrgae/qsCDKBedXqQ
aiOnMC0uytvXZO7R7+JTnZyuI69bd6dpTwLf7SYkHNjjpUvLpRxopkRvEEW2WU1C
hhm+tfpcjSoAtaKm6TFU5HvjRMJRqymlGuZlzSF48323xum9ZjUKHJgGjxuYW34m
shaqtPsqnobrBQDr/sCl1N5erkV+HbZeridpsNaemK0+cDYIiet9u3YMAq/UJVf0
IZd5GAMxHoC0N7fmK6D7q1A6MDu2vqU+iYV35spb4qDsY0Q4GdyqbvPrvS79RtBF
gfH0AfhD77BNVAkYrAP2kVMQmqG4j88LPSt78hk38XBTNuGn3u6J82213wtP3B4v
sN1pLoftroHReC9b7o+jonWQL4KVBmpqBEYhMTZHobbA+YoGknZHaQcL2QsmVffT
V9Vxa6UN0Ec3pSarqaFWg7nS29aBJdXp1FzuPs+xDDBeE8K95n46SfD9mvwqyjel
oeBFTQHZHf20pkrUocHMjNM41Y2k3dNExNaEixqHDKNFmiQpOTGK3rj0gm3Y62Ya
gdyf3EpLFKH8JMDPp5Pt9leKGDmDz2pk5PkYHFCWSdg7JcSJh/jaOlj5T6TlEciv
tnsXnTVle8Lq9NUB+lKSD94Bus/pQKqUDqFt46e7WPLqsvvxvmcVuoitUFC2cKwg
sVXqdivm3HOnsKmN8g/eR16CJYSbtOZfca+G0aNvI+9Kq3BqEh0F/Dg8TZz9uIf/
aEwkMRi7aSDUf714Gh8kuAMETbTkd97zRDc3n8/D/XmvJtDwvxVvn2GuWouVR1rP
DTMH1jOIOuCwXU/6AGu+2QAGty45w4drQadZcS1XnoA6COC7/pZ4VLgmhPF3xHoQ
Ppk1nHI4aUnfjoma/xjm9kh0C2KOlUY7sd1HRK0MLiyt/YP4Z/P5I/VTMUBYN3oG
zpS3goLoLnam6bHrQtd8nF/smSVY3d3Gw3lYXvqP+ycP8vmUX8q9V95n62LiRlWN
P9M+A4/dD3QwBbFqjX+FnUgm40hgmVOrDLEN7DPgrkYvOZ4h1MZdFfwsfLjlt2Gc
Y+cHg9iJjxfHXzqi/NCZW+226cID0iRoJ+n1K7Zd/fsIvd2hPhGmY2Vbb/Q9Cjde
VuovyHYLR2Jba2Sb122bU20OjsBqY+tRJrZ1bVDfP27JrBAMkauJadfYgknp2b9z
EKJHpaV2Hl98fmpjk7mvPsstjm08bDliI/gKRzqfMgq16fhy/Y+aPYcjqGoOcLTc
TjXLgHA9wpeGmFiGm8UXTOiSxEknNfU5VosQdUDLsJWCcopMVIwiSSK2KTm6XPc0
BzYRMmsPM4++KZyUtfa3x3lmCK7hd0ywmkjM14jFd7pcpowaXMrib7eglmeRUMyR
g+uX3tGVKOmH0YxfQJHUallTbibpmsdNfdbLrzOE3nierQwtHfXFEQY+CWeN8R/z
si4x3NtkJgldTlIXFk5BvJhvs6RqAX9bsmlLVKQ9jmV7kw7Q9mJA2mChQcHarOwn
hpQHHBXPwX7wAUgmYOfNYeX8/8G9GZ/9plwwXEeM1dbwLDdBNuvhnStqd85E70N1
u9eFdCMhWFXvo9JYeggHEGAQyUp/psWgdEj4GhdMHhXCvKlNlbutCyP3NfTk8zsF
8iSHkeuBJ06faVK1fZKinjHy8UcjhUtgKr7qnrsSbOM4upxvwHOwrPoziKtMy7Ct
cK2Qs8rtjUuSBfHqHjIkIC4hHYOv5om5Wa6T6lZ0SXTvcjVxyjkcTR58iSe03stP
vjKooJ+quZVWBSOu99MycaTK7qyyR+7QgvMstsSM5CH378xpsFEgDdnjczDJFYuw
pVlgOL6Y+Y5qfyIxu4O0IxKhE7JsmalWi1HefXbXNDWUxaoV/4bSZaHe4UeRZmGB
37B1qsj5HBB2UHjozehr0Erhy9y/zGPGIiJwS0R6yebSgH69mt+dhxhXl2adCqwD
1fsWr4JBRaB5L4j7/CoiShWanEGrL+kz+LPdokWtWjWV0JvXotioAoMklRcc6JVp
88Lau4NutH4ytiB2+Pg2KjsO+mY16k485zIDT8gb8pUB60ULOFNnnYFWNxFP4ZtQ
5N6xRnNJ5i8Deov4wB2ASfAxISoy3LOUH7WqdL+CBoZZ2hz5kT9XGy/ADubMkRaS
453CkRppsjWjERYAuzEJeIm6igIu8pVNiyASQhB6WSdXnZwFYd1rnHZrEYFQWleZ
WSgRaFPfCuJf3fdwfjLKHmWykw4Tm88Cm49tloBXVmkasWg4ZgPGcDNtG/Jwzvn+
BqhphH02rtomR0r8IktFqLRiYPwlv3tSg5bPS9a4qp54bV868ElmYEw2vUEadMr/
QHAeD5pUBIstgX+Zq/R3xZi94TWdwvC9JiruWm73yLWjcOwRYKbWkk7fenZd9rd4
zGIX9oEsZmPP0osE5UgdiD+JXLQfz+F18aZB5Ee47S8poRK/ZRit+jbvCWA7ul7E
tdvdg2jMzriV+78pduDjT9RkcNOPnrStXXUyN2B4RTqEanukrBbqKAynO1duPL+e
gwm0yRPg3wM68b0BLsCmjDv9DZ3oIdIt7OVUY4zRtQzj1SFQX9P3rgWArFHZ4Xoo
gs7+3Zb+HqEBa/epfHXi6pYTNgoIUCJY3N2Tlhhn9/lqF5IGUe6X81b4jaoFx7Lc
3g52ClkRIl2UWKjsRISsK/5On/6SiiVki5rYPPnw6DEcpgoQGLc3qwEnRLM7txr7
pWA0DroLUEQO5MXa+Msz+E3fGCFAR5tTtqA97vDk8tmg5W9XpayPtD/8KC+NSuFG
DUFIArxBWoTsZtt5XsP0GDlZhwQSfvUiq02fyYxaXa3Xg5tAaDzyRtGQFYZGk/N0
rGrASeVp0ZYJssi+p4jhEkg6llED0Ln0X2591Js5AyLjEN7/kXWZiW5mZ5xcOB1s
yUV754KiBL7SSoaNbBwpsHVuN5YsRCiQm7XXhNL4wsD0ntz31pnPcHeB7XCJHP1c
LaEr68tK0KGh81KDxrzL1kt4/SZtibqPUSXp1tupN0lKvJuZNkjXr8DlW28K9pDt
YSr3BgMjtYsAl6YqR2zq8KKyA3kWM69khDtYxwgXn7pwlcCFLs8QpgtRm6e3pfPn
dqmRQ44f58H0SzWKurVl6wjwvwjicAQ+t7Ok6Aud7+OMUQF7yoyvAzW2wSL7Hp7X
ni/3aPhuTHbpJPPDtjy6o/9DbO/QmG4eSBT4kRaJzHJaGzToPbGx8iKJPoCLWRZD
YOKBCNvT+9vKezLtrJkUcNzPJvDKMaEJ+DtONUXvDMqNBRV2rlO7zcTDMhwZqA5Z
uDwH1Vr3YjwKStrCOLxkokFdDWvAYdul0KatoVpnBQGppq/lb7b1M9WnbJunCKCQ
IRbOlzsH6Y0VdVfgDVAuNuxjcs0OMv8/cHMPmYZFUmA7WIpMzFNEcR+yBvkweypn
zmCu3Akh7Tcdzrq9Kg6jIG1LdUbStoJHJZYc7HGK6WkJco4M6yO0TprgJt/JpR+V
eMCMBedWx9b48R933tyzm2qtNBUa7WQ8lv6mZqK3eljxni9KB+3asKA6tTyqWuDt
FRtXxSHtFIyMhsQq7auBhcMD1q9X/SPCq8WRaoU2DPcqYNjPpuO4rnNf5nzSud9D
/q9zDNksoXcVnPiNmeOXUyzGEF6UcVWwGMvJBOPSD2gt0Ex2dchdR+sQZgxOBEwI
6TzExkUiOZRg8X9qasPezgPN2w7fRB0bRO3iClU69i01yF1cP0HCX4SJM3ngg0M+
l0pbrm13x87RDpeVd00zbbPlhRyYxsGDS/6oQKWuS158n6vNLjlsHcASKHSqtDfq
0P8QdeUEMhFUGzs4W3GfxHarVDOcKgQfO29PyOUC29+8B1VEGQl1PUdMkurGoQU3
oJ4YX8Kssxz0x84LdanFNS0IGw+mEgM3ccDL6kqqqlUQ15lucWYwg3vlX/QB9k5E
jg0RV9FbMmiXw3b+IqMPU4DfKwoEdbSqHutEkBZnV0VyUfTQfI2YZ2V94w+hcNut
iIzCW8tA+0QsAu4SnB4laUlT9kElUL3JVfD8cUsl7ZiXOGGu9K1wFXWe1+0DDvnf
XelNmjzgPCo4LODpz+j9aL7WBmstRJKWbZRpFFITFAAuBfeMYHwGyq/qCanKookq
PuHxiT6JD7R+ws+u/OFHP4aPKtw/NuosiQ8WBlyvSYQE1cspKOUZTLhgZLQKnmQe
7mzIaiP4sS7pg5xNPhIrS6aF/Qk5SJMGVrvjnXeXY9azjRMScNc9Wchd8EO68zXj
g0efTLX9xkuFTOzhZRkSKdmjbUITMn//6hIlYru6YoFmJQq/ToiRu7h6yRYQ4ujF
ex+MmEMDGoOk7AmTrTl6rZ2gFt3/HNp3srCsUG5560BvlMzeB2qK6mAgs3FYxKC0
rtMrzXzwNGJYchrrWdavqbjbCXfwl6tKDw8atjl8qulU0RwKWQ1n7rwBv3zPEvXS
3Dj2+DKdN3yBrpohhPAHS5esgzBW+TdpOxQ+fCJmsUYbRXahu9qoV8a1kViDrAoW
6x+1Up9BT4X85Sa/4QZ/Cvg+AHtwLhp5U6ZiJtmvmmQU8l+F5HDZazqrCHmIoXmv
jKwEZAbN9MXkRm+2F7lMbMNYht6l4kZFVEYP/601HZ6fzaRJzydnVDNj2a9d7Apk
Ze7wqJ7z/1KVkMMdkjV7UsaHAAdSAvRNM/TtONUhQrKTVPiZp8F9UYgOQV/iFRsU
RtnsrUAgniFtGX97hx49HPBoMWqVybiaYZ9srtRTi4lzHsTsJ41wvSawuFAFcHAN
Dgx6Ll24g3ZZwQEeMJuKC/otSR5iuGrZdFYzEKCFipLUiKnQWV91N5J03n4glnDR
3xZY29iuQVFtiR9Ac2WetLXrKPhKk6sq6j1lyIysAALuXpg+06gaLw7xgi0s+22x
DFLOEYleyJw1Lbf0M/+zIGxX/db8M48RV3wLpVfylJgyykI2BfFqJA9bg/7c/dP3
dp4IBhOe0LmRlDKOOnesVSPjpVxW8BKnNxOEdYKvsETN/lddCSYq3i+ufN+C91fv
RzNDcBHOwQj4X6Nbk0UpokMIiiv46oCLmTalRCMoR/NifRa9p3XbIe6rKd2pOrvB
CKc4bkQI62Z37fRy3Gi+RI2mKljUQZEes4Hhq8hEsr5O7lHCUc4Y66s0itV8Qpjs
VhtjWi1+0gvF1Tb7u97KGppivEfMaKc/jf3XPFYXolJHGh56pTvwpLa1tXkzjgSM
+yocduQk4L0ByY6Durp+nT9VyJrLprD11nNBOLZd0EHuNzmvAT2WObr0dQqZR43m
KsAmg34Gj3GfEbYkylKT2Qb5XtyYbhhRffDPEGmiYyAHXSAbUPYlSBhgN7UAK2UE
44LgWm9Ek/AkssTiOHjLUolP3YRG+I+QSwD40DbdYwzf9YLfKrliwI899bcuTMro
6onZgMWU1+NbUBt5jvZwYCD9dtMqZicmMXeb8KnM1Ii5eHYNQ8bpWCMjudiFZEJW
zcYdko0E4LE3DlPUiIpZ5VlH/TZX6gVC2ffwqT4vb2SA6hyiSLxT3bhbMxb0og5W
51NgA3x84GrEOS7m4A0IoEjJz1D1pKVp1GOraqFFhRhTDWp85Ourx1zo9Q2yeNYe
N/NWZVDasMACUQ5DEfVdsj+IrfmZvKhr31Tz25oraAcNMFT+8D2L3gWTS0fOlGqu
awNO43PNSc8DIMoYqcXMw3/WZ6TpuDWPVKg8ABq9qGdYhNjT0gqFj7DtP5GG3uXT
JVNy+x2juBx5doPBT8ns/8kAAJ0PxsB6RvU+UuOoyoG19LvI7X9KWq6AC6y4KiPM
JIv2xwegzWEqogS/y8MDyXxE0Qo+ZjpZQJp+ss2jveqRbi+5smC5TrARVbpF/x8w
hChwqgLu1pFbxVdYxziHDSlBTgI9DiKHwKPqrijGaeU5oKdCh4djPjYyvbh87KaO
K/fn8xP0eWtD58wb1EiH5LQAzIxIHb8M51grtp8OJjK0gLR3dPgcFqSzi/zGQSMH
B1tqVslAKOE1KINSy9IDf6MNhIknNuKNpBe3WLEDwHu0RIzPCsaAc1mJkdUNT3cJ
eJbeHZo+3LerxsmquUIK/7PDVkdekFK4RNdO+srF34+4C7q/TcvqcKcFWP4aYe0p
1w4fVAYnvQuqbNAAjAanKlbKrZT0giWDC+iQOuSnDXuF1pq9WrnPPJp89A6v7SCZ
axDbRqvFUBfjINrr40kWWgovokBUI+Ccfh6r53s2kCSKrPs8XrrFCnfUMYaxRK5m
dpk7dL/J0tG0JIJEp++86BMgiWbF3n3MWoF5fiuIrWleMoGHD/vGYa4a8+pl/01L
yuQHf0zeyGcmFEbWCIKKIwkgd3g4sq7n00Cm59DnPiI8ywD/uD9aDVSW1STj0ats
F7mOqttrHg04KO88ODLrjrbikfbTjinKNFetYts16xJoEkCL3Em8q/EITK1y97NC
EmK1qqZB/FsUvKNFbj9AIH6poXhnvzY0Zppb8NzELdMAXLW0bawEQ8WGFUfjViFU
IMNRsD69uDCVHeQQt9hNHS9eLwaYVvQJqCMLBKrxBohzAhQpl+T2EfJO0836NIiD
H+Iq2UEWlqBWjgLNLHMakSrZv+zqVuVueA0KalL/UKQbjTW3v9k7qRK+lovlBYPc
zlfwgqMnGZS5bJZpX3sxj4dQq/sbsmt6IDgk74Rt+ZlbKbQCeK2Nnyz6yNY9FUOL
Bi5Ug2rgMCNPpDOX7iLxso2QnDzw6V/O6B3YCUFwa2JYl96bCzRvy5JKbKT4dFIA
ag/FbOowzLWROntvuiep7EUT2GHYd6le+lyAlZgvwuTWOMn9ZuZE0fi7Q0VCEwFU
VxErIJP2uJYE2Cjcy9/37Kg4pO5MPdMEs7TjMFL+DPs3F+tGfiNrMEkh9KFqgpau
BX9s32cgkC9YhB/NN7CBWw0hgG1Dftd0qrSHGGvXFLu18ktGMTm5/dFxfdXLWwpk
JkUl0+7VKo4vHyojonW4TbaHtXNKaXif0SD4bSMQ5JJfKtPmb9hur7sXGJzyVq6B
lxJFWyUGFRtOC44GeA5pBM4YOfTPF+crbv2WMQ4ZXkqtHQcCJSU0gM39pNYlXqJC
6+4UBG4BhNAbmmXwDSraRdb6Z/hAko72sk8H/RRgdpn6uiuZBC87tgz7Z5c6H9vJ
yKzW10WMQC4R9evj5ReAAtVmZRBaiMcAfYQRsqIUGAWkQ/qTWe8nbbEBYouJcvEr
RLBpeYhmO4ND3G7W2fkAvvgkpIvcRMfPXq4nyjdOH9DxkmB6j5vcvnYsi11ogrO3
Zwt1fiGTyEP88beM2pCiflFBuH2LOpRbGXR2fNStUt/dEf51fys2IMSejefviqf+
fjMOD1p2SFasRy0/shlqFxy3FlAp+y9t+Yus0rRTEZhMc+Viw8Lj6IiAC4A2UUi/
H2TP4rp4iXL+/NqLvJkq1CQ94VgtkPz8WIwZuL/WxI/Pr5UVPpK9ucIUaebken5v
M/snNewgfD+aeX8eUYRG6LtAq42XfDyNxKL5nkW0IGUfCLcp0gH4tU/ZTlZEpyeM
trG2NtoOzmmXIbeREVd+9FgLdZqg21+/d7ynVbK83TEfFVaXWgEX6N6ZYbXIl74u
oWgs2L+hWbMkk2hvr8G96oGtaPDTslMSQjFkdOHA0viEZXsWWXqrUcHbAWTpNoj4
d9pkC3XDsqj2Z0hcCLhRMQ9IP8vIrBHSGbf56MGLKzbmW97dA23Q77/rxITb+d5w
Lt8uqzzRCCDWgV5U5d9tcASZEw0DBLUNs/90D7P24LDzkJMuTgcF7Tt2A0OJ/QZ/
IiOKB5xoGQqyWWxSzXkupI/WIAON93KbYqxV3pFxV50EsrEDVP50wHB9RbfsAJ8r
bT2gz+oiH4AOjhj5AWkmXAnDFXMZokBwvWpiAYVLW3b1IKCI7n94jCQsmVZAjKd/
85/2FD+zK+WobvFG1T+y5jaQB8lLpV+prTjuBCkG5MYKOyGV2qequUmwGUuZVsUx
Qqihw1Ft9I8lmvHkdgmztcrMjVddwP/VXGUZPrOnRf4qfYroY/lsyatN/OUkwWkR
Nj44Kh3/+Ndp0/z10hH+bzeFYHEfUfSP0S3JZeiGQHQndcpck9qqA77+8lzebxQa
NRPfePB4YbOCEBeQRyQIc79uDmkjhtnqLRXnu0+cXIZ0FVAFQ6MpYBhyocW4eWBq
ol7s5aGwyT/J3HtPvRGRahcQliUmR4jskoT5Lk088Q+eG3G9NiMz3U1MsPDPUcah
TGdY3a8GiehQet14WmGcWraGMw6XxAP+Y17kRQejFdDmldVLE/eY920ESSBrzJkN
GGZUCwUdzP93xz5pwgPxURipTUA08gdKlscNTI1/ULmITOWYf0Nb5IshRv2fGCOf
ry1DNE3WHezaoQ1dPPCtnOG0ShcO5WH2i7aAbRaiUVdFqNSN9w0LXOSOC5Pex4iE
zbnTefxfc+6SZ0Nz1BdxRdI2aBFJrK9RgmpUMM0YUB84Qsjo/zr0c+2YKwCflsPZ
mXSKNFLnJ95Ogp1XR+uhlvIflpQsSm31oh2XTEJ+4IQMIrshx+ep2azg8wJf4qGh
8KA8fPM3Vl5O7YZtYUKXu9PT+JWGsEG+5/bWScLaaScdR7W4bNj4MqxvX1XGnhDB
pSJQV8xMpFi59B4l75U6EVB/z5nIZv+L0EDdjK7tS5eJGQeNGPUBQuxDsBxnAM6R
jgf+UzYfcaUmIyn6I4xst4Ykh8aJMUkFhIPoiZQi3Yxg5VhiYdS1WAU4rn4FX7e4
HT4EdzBrZ3TyC7I3TlaIkRaq+HVCcqseWRVxfc8viNVzqpXgyOPKMeACAp4i76cs
VT2sYxFexScryw6H9S0X35a5e9vbKy4L99lDkBC+jyRWpkQoyYlXKig2j9AYAMBM
YUfuIVNiDNeNJ4/XdKpU6ppiapPUXPHdicoW+o+AHZM6uQeqxfG4Fs3WOz02ymJP
4oBzkBmEeuPw8rIkHqNUfMmIeo/HJyoTeaZjJM6W8Jd8Qup5JqHCk/0r99hlsvRW
15KvQ7bn+T93IS0mBzY1t3bNlgZJKenFKhGyeVg058zbVli5VEqjw7+XWADnSiR7
GZWlq9FXKefhHOQrjZJyXoKziHwe/2/vN+Wi+8c5f27WDaq2fR7iPueYsw4VSge+
gfnfQcLrGO7V2702H8mSOxiVUBsQJWFM8Jk15AMCit+L0JNU32y5QYLJyrU5aYr4
eP4A6BFt2q6pZhwbGB2KLLK/su2o0GXTbVlGDHNG5zOERKHoqYZGC3No/60fF4jU
bcW4nyob97MI5KniCGsD635mKCNgvxihKef138xSNFqQY9mRTqMv2dhVdOgpTtsJ
7YOMZhmpEazynKTr6vAFPGTtxUAHVoz2mwTAHjCpd4CWmif9MbF6/8GuOzOEj5BD
FyZBxfBwJr5e0u2cWCip1SjWblU5eqUJh3kr1lIN3TElSKFt8zYaQPlHgeLIX1qD
+ZwAIFhe8UamRTM1wGXDbOO84+nUozQsVbZssK0kz0wa5EgzzyElBopGeaunmOv2
EneE24/9HFn8PjL+Tf8Nvegyv4tdrs9wB0QcYonDrnuaEJub/zMkBA32V5YrlhgG
PHTRlGl8AisAuYFuOkfSSwn6dWXORRGBBAed4W6dMmPwG9WLPp4sZO7LvDZLTc+T
6VCOvOEhH1aHTA8mkESTKIgKEiqaqMJth4ldm+O4bQ+Me1SDRutSdRusEeLcmzgB
fyIYtrMDIw/rkePlsN4fnI+59cenGMYZdI1Sdd8wLScvTWZl9L9Gwgq9weP7FECL
XvNgBGV6WOgpXkBYL/M3Hq3CxfCQeD5xTUaGpoeeHhaAJZ/15sdXPYXCleCOKD2f
USn6Wdm/r138ZKEpeS6YgWSEpeVIbeIxGw6+ap14QrfobOqlNU9QWcUpieHl0lNL
qYs3GwOaQ+t8mHn73NwGNHSSISYB8q2QjDDeMUAqvDzFUPyofmgUUaVssy0qLa6u
4qxVdU7seu7rvyO9CkzchcCXHuE8B0bQ8eBZioRJriAm8aJSzFhYeqVQFQo3J7/w
NGQZYtzTN669hkIRwDtPQKfiK8Q6/NsQAHjt8pKPElop1IoE+yHFxDeWU6M6Ax6n
vKmHcor8TE2myZWlWpdmRtyRzgNFGvogWIdyOtcoEnm3IySqHB0YzUafaizCV8Yg
P0PyMYZp2RJJsfQiT2WBIBAf5NR5l1mOXjPHchDMF1iQdVGu6lEvAG7OU6YiujTL
kNdtFQPlKsuygn9IP0sf3m5v6/U0T/1jMQwyd5O4knsR7YolqZJLncwJXVhDad1Q
QuKJUB+e6/iUHLHAOZr8Q8W5cPsPMbhpkm8EgQmJLfTwtwNfgebVN3rU8mx3Ih1N
Uw9PAfbyy2vAqTHvEwiS3HTbvgJI6ULfXuRnhlBAnPvnSajq7S6c8yYMrXoVVrKq
/2JI0G1btDHQ+bFbiEa7bfkUuAWPeMmsYkyl/7iCsXj5GA+NFKV7k4Jg1gpHhhqU
ELelAmNbOwkcT1gbv4KXzpokRPSmZkpXrySWCAoU9phj+GcmCxVNPWfZUfwIO+LQ
FhgLogD9w1PEmADcKhaSyMQVAD8lykgEV6E/SfRPQsLeoPW/uQ3ZsPzQHcJJWV4N
c0wWc7FQAKQ13eGUvmjWdELayMvxV7XdIOPMjeyXIspvduoOBHoTrVXKeJL58bJQ
XieB8XmkusEqQQJyO6j6FhgHJn/cjpoT9aEK3leQVB4gyUYDIGhPsVAgbkTC1bSf
FXHIYDnhie/xwqbLa5tJO8S8bvsEIwR7RBNY+bgbtVDyYgDbe8TTBR/HfBHTivGa
EbLaGQL63mOnyi/6fGN7KT40/k74BIyyxB41yNYzkofYXYWjmxoBZ4D8XtKSbjmT
0feI23CAsZmdfLm5PxcfMTkIgnzPSo1hyautvo/QO1yB4m36l49fI6lbwzaJi2nq
97OCCg5/EqsQS8r0aM0rXkFxMZ7fonrLS/Dbt0jHPbKFlQZ2YCD/2XffCe11uQB3
AgdPUHVrLJUCkcVbUMt0ovR1Zk/GU5273vivQbQE56rT5+ZCrmqzYE+4B1qQi2FO
N7JKXIENiRVKMKEOs5r1RJ1pZf98gUvr2s7a6z2XI0l8WcQgKm9DtzYDSymSu6xa
YVnwIu8Q1+13EsU5Z5N4UwdrC2oFjRmzBZXOzhAVf7RY73YvJ520lN7MZdVIlujL
2PHhUfCnn1ZiJMRDhx/OnQ8kfx9lubk9pRlhNH3BAZkwjKDBhD62LgTBRYgM4txt
vbgK2BvX48HfPonY1rke42IH5EfAJyOibWLGhbdyEKIEkqIQcRu+N9Y54gkU4oVQ
UR8w8p/mYltJoEnUL9tkKG8i4FgxtN6p1iwJpf1OYjUxeUPGSRQQyxMpFS3qba1u
c3KWzVKtnebbdgRsr1vk30ky4/PnM8ZO9KKPkEhvVxgy1raadqJ/8hZihLXBVtE3
zbCU1hUIMsqCCi6EQ/o4ViyLzdt8Ybb7TMXSGL9KJxhpoTWgz/oMzv7yeNqKoMXG
bKb6SIkiW12BorG9D5W0lHANUzOO4Jc4HIw88+PcnumNfNa0z5x2i1nIDClQATeo
25vNhIBnaJfNQKZdO8Y/FV+9GpxI3Mtgmb92/W48tJIOU2Pjb/W+aMHicuJwlUIB
LsRKWNnRKOLtypD3/0Vs8zzrHu0lynaxC7peHH9GsOOKHBNzB5wDjwtSLfDKp2Wt
icxqYpS+OMuKFZJ+lgw4wZH2rEmz7bsH/S3uNg4XWRkBJl3e3zG2ykiSrmcelKKn
Q3+R3G6oC2sK3bIMOSkqwtSv6rgIqH1I9dYmPjKSTtsAvqiTT4fpUr7v5wgF7Adr
nutOSu3CCyLToykf82KlQcdepf9FXgxQAyrE73duaPQw0nMSJlh+4ddZ0RvdRUDE
ZpP0WGLGyxj7+1Or0sNua7SnPNnY4ineGKTFIaJPXj2K2WRw1oTzlJOZmE+aVL7j
fBBaO45z+03rnQjrYAqYX779UdFH6yyDl6YYneHUfazQRqb+9Gw4Ug8fTTvHtANc
A/qOqe6qyi3YsBYbNuaQlCkwtiVGahEtqD3AZucxtqP+R8pJjzIdKlxpxS//Mkfu
OiyYWN6pGVh5Lfl+iQG9Y2Jww5a2GgHUgdt0m6GmsQRfX6DvH1P5mE4zE/Cu7HwD
HjW0/NaV9NmlwHrxYU3s6KTkmLlsADK+0TtDayVHFgmhDKlaZot91oJPmQMLgvzF
TcyezBFqP+v3ZpZZ0/X7LaMhPd0SLz+Yhj4O1a4zvyZBmno7Jp6wfmFu4di+GlL1
82+B4+DPq8SAb1QmbyY4NWzTysygmxCkYVAHgBMlMR3lWWyqIKIEU9ev3p5jAcBu
hqo6G/bdluiDwYg/x+FuHZKATdVfiCnkMwmvlqixEqlzrfzqJXd6YPwRvwF7BeKk
F4yOqHRvKvUCXM/H1bRn536IYBWwOSMvgx6U9B96nOLAzCeUcfaq3JacKZ5UcM2w
ELM4+ppJTYcQGD0zJ9eIaHzXZsU1mvdiMcFCUWo57bzgvYtQVXnJ5MnvXR82rGeC
hBPH2t2rrUVlkOEfX/cjeDIV5cf3ZuMQcSYKOHrOeQgLFEIBUqY5VsqcnzHOMaPA
jZZBW6n2fASpnkHqDf+DIc1fnPpVbR1XbPxJAYe1Tc7LWPpu3cZNRuGTtvDbfOcS
3UvGgThb8QO1xmwjKtfQrt6c4HwOYBQGDxhFx8HURXX8H12T+C6kb2NjSzXEQmC5
ND/8uaUbx7RkEVhdO3gt4+BSeYX5/GsUCVTW4lOR0nZHwVZ/mOJr5i7KsXaMD7Eb
PWtMSGAD1CYKqkDI45B88ugXchkxPsikyvMlapimhH4D4Q3Z8h4+hUS3R72NugVS
D8TUWkJrDm7QwR5y95IoH5MXNgxLbCPMHJEvXZpP9LMbqkPxGt+xGj5gjRiDA+5o
wsunZXf8uBaUClgGI7LSxIhyCDGl/fU32a7hdNE+92IMWgbU1T0PqtxSRJ5VXdlN
eNiT+8bZoSjdnCxopKjICmCO35GsGItIU8fs+vFv/uvMH7Qlw01TW4Ni5TzeN6JU
oliSzOeDbEYJNtMnG5fm+2GgX5o9FI6TFcsUKImQY+knvoUQifYgkYACLECu1RmS
lTm7QWRpuRPZchZlDSEmdXSxVdZ8j7s/1Qup8gfz0OuqRm5sST1KBZetp5MyOCdR
W8+4/T7+426qAj8jNAswVeF+8bQJdK2SY/XaSndVk7BSNiw1kk/QQlWFj6K2Zw2q
nI775Qfpn+pqx3EzIdcNRTMQUZ2dJP1QDjZCAuzUTWvRYjHYe99QycZsJQEUQmom
arPFkgahJGtL7B/L85cswE2gr5R+AumMOtf/790WJEtV7YFk5iCeNb4qFIFifoUa
3bQSmWGTeCDklxzAFwOIoeIgi+iWALT44pccspzX1h5225OcuoWWdps+tu+jlvE3
FakxPkF8vTQ6F6jDfx+HQwhBCN/o+SvBMy+fwJCfFmgP4C2tzPRtU3/FNpvKJdFR
auVKvwg947b+NPdnVFAudhw2lrHuiWnGGNAoGn3PTXKDIIrDyBW+xBHelf67xNAH
4nHMwGtRJQw2+DfRJmySxZqJTWtg5CXQuwEOp3qFrjvzj8naqukD2+NGwgOi6B3A
MToAWLj05SJ3rqSSeF2opJS13TSAj+yv76Jshdo4o/Qr9+34vSthpNAkp7LxnaVv
ivT5isFeNSkg4fBV7eM3CkdHDmRUJqn0I26gOTxdnvzC6MvqjceU43R1sCywMDj/
QjYMZ3Ai8r+hP2UbBH4yn57tv5pIsBRm44HRVg81Yj6eMmyMYDHeKiA0kqTzrUNp
6bi1e1K6zlRBu/cbGBXneCovuCtBT39ejtCNLBeaZRSDskAyNb+3CFtnURQ1vsoJ
WFgCrtHRF5Dy1DxasOcrgLwTyR7vfpI42akOvdU9vB1kXvB9DL5sg2udO+LjQPvA
jvQVRScZlruETqC7+noxpjQYCPDzaeyteP4u4Z4uIfWDqTA1DJGwBDDghn7C9bXE
vUuUUSz/W9TSYMG+VojpgaORpt+4nc4J56ZNMQ8EfKdvRivTI+Qnq8IFxSPQ3AEh
ov8ZSBqNNz4FoCl0JVVaR9IWcONNVvtx5Y1zvOc32EoIkNQPjQ2uSyg2R/d3pPHN
dggfZko8zf96Z2QR5bhE7Vve2HT2Bi/s7D0WHsRH24HueIoBIshTgwS9A6tZ8RO5
U8YyBZM3K2sepeMFuB1FnIymCK6HDY4ivWdeq3owOmkfoPdNPYMO4uxe+WhWBV1O
jj9TTxB6OFWYZRcHM4vrCoGLLZy9geztSLxfGgZ0CHGUmUMDaeDEqWoe8qYDhYVt
gz47h36PoAR9BWkc7tAIeBXFX+1C+YAyNWAvmLPG2KzzimIE8MaLkWGi3SlNhhGJ
yIzyQtXbIvk+djMw/IuAn0HE+HvY6WCyT1i4n5g3mdnhMqRyILuSMPoU2FPw6rXu
jS90s2PVsW6dyPG87V58GDT1PQynMnwTLHpeMXMtYrUUl8Xta5Rjbh4v8cH6dWHI
ingGQ/FE4H8pqguipsyOsdTeCt/JAnNzhb7exLZo245jDsM0K+mzYZ1GMDseJP3t
/t6DbA3U+bBBMBusMooFKg9YpMO8TU7zekzjMN36YZo3ZUaQ1RMEZOO5IhmIwAb5
ConkJGlTARP+3r0PCeEvnAUJgzCoKr9vtYvZFBQxd4Dx84zOUZu27uANKv5y4jep
KL7LydDA8JBpRKTdPHLLsRKsPEdx8oVjBILzKZhwgCPNPkTv7M0Hd7W0gZpfosbd
n8skw5Ey+uQV57e4fEEHIDnUusMh8XCCR3mgyg0kpU7MuoX8XX+73fHknaY/HbXw
A3VrmwvRoFkqdHj2L0hcRUNHrXL3Jy2SHa8hvVwrD68EFlQ8XXWs+Y5A4I895ZqE
vR9AQx+E/2vAwA10ctznHsBTQ1fHFJkX064wdWnUmZkaO/V7ZeU5W+Ut9GikoRQJ
XDb0JK76lP0KorAh8nKjvpDbPZdTqfP0CXR8/2VMPGBn8+WqZzm/8yDGZeIZjtCE
j6NWKfjmx6fjrDxzWb2MHbvnlp4D5tAg2yQTISyz+2uSJeo/pR1TbyudIMot6LLg
lIT6iKQkHwaNOcjkUR7stiS3392gOuEHWCc+4f7bspvP4aE1XTM1oAJSoc1rbe9o
Ygz0SNzMrcuSLIUT76pc3FFIIM+oqUvMseFBH+YLz0V3DWv99CiqZ0IeZjLv954Y
fUpwKKr64LGzko1S1VDUBYRKpmWGzjx1NRwAS9H6Wb96Ln3lehRpzCXuZLVn0u5N
Wj3B+q7nHQOLFovLeXpmPVjcdj7dwWGlkVbcVENKuDXFyFF/89Xe6gBXDdXxlUMu
g6dpdhRAx5BNgDtVcVAuB3iHG/yC/ACLBWeWn7aBZFXk5rURHLIPjMF+aDdjBkAq
/E3iRN93DWUnC6SANADjMsdCldAotzsgvPg+YROlfpDQO+WDmIgJ3SNtZw9wISOi
D6Aid4pjkW5VbH9GGSlZp/jRraQ/CeYEyv3mg8sNurJ8WbS4ehPlkO5ExDZo2U0W
zqcasQbqc8x5xWjyfuS1NhHUrlGi41Cdc2RY4m0TW49xU7BU+apYsa4yWCmDQtOp
milVvd18xqmEYmz+pnKqFTYPpdQAyY9/Mg5eMfQ3qWloNZ7xRcmpb1hhgdrGnW7F
sNKZyuJZdAY7YUb05E0b5DTBRaksiD0Hfw9z8DjTdrOmcEbwriRAaAno7gWaLahz
iBqgBnnpgMNkcOWULOiuHSX+QmMXo1wMBl1O6n6HUVJAiSicdxlQ2jAc6cwtLPBE
tBu3VVWabjxD3aJKiNaK5SR+6/HeX+J1BRcBD3ICT+eXOH+YuGiKOrknJevUWAGZ
+Kw3CDCstxvd9TelELZl+gbQ+2uVfsEl2pdEmoB/TmLHRTBI3IzlF5FRIdZ+3bt+
GhlEA3tVu7I/rFq9boqIeXy1UkzqyIqt//u8EPrDxGuy0iLS00r/lSZIRRSWBoLU
CwvDgtZ858UuuoJdROOTHcs/bn05o97XgYSY6c0f1QYf5/supcRxYnNzn+DG+x5w
PmUFPWloH9WAmaa/MYzIuh2aDVq+1aiG56EGJ5SHuNIzI95jKcwO8w3UQ1HnxQhM
FMRZrDQQ2Y/9rSsp/6EfOhWwqdcuCzmUX3zOE/SbCBlNZE/h82JdmyCWbt65YOlW
3ncOo4IeoD47FjldEeuH8KYPZhF520fHb4db/kuDs3t3lVvWB1/XL6EBMBFfxYHL
+z1R7SHu2XbfmF244LX0aKXr6N+foIu7Ay1x9BalgTWkhg3ZhLt41LCSCyq5YlTe
ecamDk4ZFrQyI8KbAG6JhdN6OhysXWpfrd5yOGPmaOP4twEjIg9oSYl0InArb3B/
IDbbF6N/KrZirRxr0+s0jQMz9tQUzhzAfzkstt8jApRSqyx/hoT8x/Kh1REBp49u
JIy0/B5oCN+taqll7f0jppkepZ+LUTQyAD1Svdbj87i0Cihhd0n1Vag9vExE5VWm
3U9rHB0VoBCfNYD7ms4D4JFaHxZTmUF7iWiA1HbPdMrTfxSPqKIGn9OJicJZRAiz
fmLagDi5yd9Ly1YzPgM/B0iQBloEswkZi9EuBTD+sEbDvr58UnLBIEYIQg3csD2x
+JVJzxw1M7AQhz/OcICLqBenBV3ENv+wPt05JM/Vd619qytdr8WB+uaUfhy6skpx
ozmD/Z2P096RRnQk8dKpNxtMD+Z6BfyJLxti+Dy4qUjsjFRyp7+btm4fupJ3vZLM
1Ru/9jAxycqCoNxcsrd8woA81JehuKheUF/AlPv33AuZKCntqS8PqZLUT+YUjUZQ
VABD+2drf0Oz6JSO0uFckQ4YXtqEJjEGZGV1nz+zqw5e/ZL2xeUBarluzuaOOekD
6dqQmDIFhngCsotduRJ3dhViTuK9YSui6MQgszVQOpPFu+wJBRsVmIj0noSkq469
WHiadz4dbJZEGte3EJHv+tuDlAVLBYZnLgDeiZqsW3weK0c9JE5nDbkGz3rf8ukw
yicx1Fq6jViYZbwN8oO52XWRaVhfzkg5M54Qf3wd9X3Q87GJrXCqwHkXTVzy8qbR
kVA69urNAh1X+TzY3uJM45NMT22goDbljB2LWl/jlGMg6GvSb05IuxeWYWPAPCst
J+ZqXynyNNvZPSg8vXrg21REx7F83eBXmJANT6CuPLfYpiedjcSAvTiJarQ857//
e60aPJ6gvga/J6Qda7ZYLEHFcAcR0meKsuXl31pp/0ffuBwfK6k4h+ZTFPgGmiVQ
w5GlbCl7N/kajHa1tFeenlmDvmxSDKH1fcPY1srd1Wgv9IZeBZV2tCS6gGFgMXSI
/ZsImvNQ3aV4ECqIW65SUWzrhZt2XAyMyZUmM3lI/l8NJVn7z6gxDnQPJcKelU0E
HTjSs31BuU3E8v2pBBURQYClfTpbQ29YzfRgjzQLxkVxV09PUA62LJXSpUXyCnBY
RBm1EUWucmw+WdJCxOahOhwfyTEKxtn/Vri/KGgbURv4BpPVBkWUiArC4R+rDwNb
UE28D9X66cVXpkg0etjr0/wugtsd+TwROx+JE/QHSa1FlgVwh7ZxAUjLPYCcF2dd
qt0h3edYYlqfu+/MhlaTKD9kruQg6eTywO5d7uthgiVriYixG/LuxVYGpquVWBeY
QtTBDuYlEACY0XfLggzmaqvXmYzA/+rBNpGY2z2+VGjAk0j4JruAFTAvExCIFaS0
Ky1WSAOCGP6Z71CFjS8bfQZ+Mm9rIvhelSIXVHx5v7qXDCkPhoL/B4csctKVMYoC
eqsNwOj1zj5smxG/s6FA7qszTMW7suTtBfQPxwRfZnmbftnuvFrLWpzV6t9S+Gi2
Sg6fhHkEpQ11bRHmaezpF+toU7GhCwP4ebeXSb6ucNiW5TxgH8cjbnz9x2zeprgT
vHHwdQHy0hAbAta4DBmIj44P35yovRd7lpzmhTxe4AJkzbqQUwl4ayopRIkpyRUa
Kb+ycYgtyR7poWvrfcUysPxZGsvmHWC5PsNiQ+djNXJhk6dMrPYUAjhjnrsjGQj3
fNCJKL3drwHOYZbWqQQ1MiEacA6lt5YNPV7yVC/1LBXNKydYuw+gEp+emt54vs7s
pBaQBA3z5gYIyk6PYe5bc//pDyayNV01DEt/JcAmKtBIJCQsYe0gjExv8mnfqtfm
iOfbah9mJT0ceCcPQgCf8CbYTiJzBG1J8Qw/H+rdyJ4Lhg1j5YCkCpRmSr566rk4
qODmry8PyfcVc2IEd6sT0dvZx5WYRwAjssJtYicswrqLU0OgjlJhnc0k7dQDPtLq
CcoU9fICVmKcfK2HwF9eNuPBl4r3hYGCqF3Tb4wdGQrwftT42Fi7uSjtFeo9v9bj
tKW2MLm+Ek6NFTtb5MvW/CbSIV5b8HJluk0pKe4ZjZZWLBPtdo+vq6bueo4t61dp
xzvT6sqg968JNgbxS22NwvMGFuZ4gaWqXRIbWxYx4a6TT0gTo6wBWVJAz7xvsKMt
5nMh+eRTcOB6slSpXmZ6zNZkI+24iJT/Mc51QrYV/CiL+VGOvHO6mmkBp6ZZ9Wnx
ZpjwLqzEMkJACnKEMXdibKL94VTS1Mbxs/ulJVVZ8zJzKri9uQDP6W04B89PsBrt
AQauimcdlTZWp00TzgdCRLCnG4w5q3Bblw1r8P4cpsNIq1pNIKIDP4RFEzh5vcxC
XF5FTxSqOuiTwT3udtRJ6ecNEw2tpAZeBWBE7/H6ZADCgHbIoTfmGo0Y6Q62DUuf
/n6Z6VvTEs1B9s7Sy4PjN4T2NfZ0qY26BCxWBBHOZC+1LUDh4V9WyHOkTK1oJcsn
E6KFSI70aPOn2TVL329yVxX+V+NQWLzDVdhEoa9gvojS5hv0E0FU615gLET1WVwQ
ydsP0ZOF+IQNs48ZL+EP7Onhst7OM/1199v1SfDsFxs7dtga7yCPIb3OewsjOAPz
N8wnwLmNvEh9TjR2RzHoR24ILXl9hKhNEkiZ9nfb6fU+BBybiT5nbwdreSCegJKn
4ohyRuQWFLmfxY7COQIY0bKjWXPjMAuvQAMjgR9fIfinU5M3lbxsrbX7mzgs0bF6
bneNLNiYQmWYQC0x+nXzZnoHmL5ffOR8M0tfVXPHRf9OHzcxL7nRHtqunm6IA0JE
7RQBsmdMMVSeXZE/Oz5p6iEUkl8apD2xGFMZCf3V4Qp7dDTFSg1d7KnHXWzRB0TL
/fPuMSiJPFhrBM3bGauacNndGhYeSw2CHkCLhRXDXK+AIcVGmDTAoVLDiSRzVEKF
EigWE7emEfM2y+RMvfcuCdBK2ltWsIeT/9QjLTCKMm3Ozp7mR0kQ1cwkFvG8F0u0
w8V/XTEwcpHXmoIsjBIdITC/E15PTjfjY3UL29xRgtRSj0U9RWoH6wkUUZNdbO8h
d70kCdPJOlrOrbcfVc9OiLbX7w9MfDM7Obyqyln8TjrDnjHzTE5EQ7XkEmt0JKkp
32dyrVB8qzbCnyT+GtHOIJA+H2kPmovs7KziOF5BdcRl/XyMh8UhiQOBW6NmBGwo
1IEkuIn+ydgbhqQcyIlwU4FFoG1+Z/rghvQ1+kEYFdRidkF9yah0hadl00tNIufg
eQFRg77eXUsVCytGXe2mF2u/Aj1O9ZUrw0wRB9pwk1UCBHqBlCVjHz1xW9ukYFSU
7qv9LuPk3als+Sq1DCEclxz9A1IhWn4ClupZJxaSUoTBGJ17iPZ1DeibWtrVBcGR
idAAzJgKwz2brGy/hDOvuVBelPcHIeTXkhtt5sOcikyBHrBcotmjSrmd57vOe6ME
q3BNZMYN4cDlg5lOuAH24hOD5PNErgxX8kYoKS1XfxJ+kJTzO6OQqNI4o61/+Yqd
Vy6Enc+j5GLDCpOFLgWgMqkJUaSxQIikcaJowwHEVscDxb3BeTn4McVLQshzWvXP
fXSwhtEJgKiFgCgTIRdSSRJOdX5LZvZqjjnKI1/5qwe+5zxkU9ZiwbsD/icVHB0s
P3lR894FKqc6qKID2O5tAPCb55NAS5sG7dv0+sCNhGmPLnBQRRyHShDzw5jAPPQA
p0NhFAPUGCuRFO0zsSqDMnlyFsfjc2odLWpyAaoCb49aurxTWkP8s7FFvyyv/6B8
WYJkF5C/Zu6idiTppufoQjCD0eKAQQnBQcjCSu4S6FCiN9xAg0bVZiJjT9tRH9XF
xNjEzCR+YgGBhrlNlfbQAb152O2MrY+zUt8MpEAd9zPKzUyxXMR+FcCvEhchWIRe
ep5QY5mptxyA7SqrdHyZvjnpi2l26BQamgi+TVQE5Z+NGsOZxE3VNfT/5xILkM3p
Z306qwJB3nijlXjRaZLnluGUI9dZIQQGSNZ45TO2jPtBy65SsFgz4+Ro4/ISYMOw
Dgf5Tym2eYZnbfsYtvkZ2yXGbIavjxk6nOhgHNzbPudiX2JUGYpn11/lF94+jwAZ
fMOjMyo/ipZf5eTaJcDhsVDyzH6qx+SyY15eJbOPm8dxJd23YL9bzxDFrqXaFAiW
GYc7s29D9HLhh6hiolWzgm1TIocWZFD+q7YtVgOSleHCAjs1iDaeVYd9T0g7sQP6
OGV1GcLMl1bihPFjURdasXULcwTpN7HUTRQlYp+Baic1eSRu2L/AdUSH2BUt+tQ/
8DjwklVRxKg3chhW3+XyK9zaKNh1vwdxMPiJzov7F45USXU+zrHB+FriIOYTlj16
uVEjBkPRZ98XAeSTCPeUECuiTH8otUqLaSVubLI2l5o+OckKDVpdG6onOuW1Bcw4
jyuDA7KDSEizlBax6m8ZhcD9tmTU4KUJ0ZHA2wM79W5OTs7a9Lsam1doyh/uiVWO
u+diDKIheEEbHDUq2E2cIlT9LPb+mAAxW/OxuXCjF7DNbQDzDJ6BIoSzr1zY0EEP
CoZjLWmUlAti/F9umsEZIkkA4Tsgpy+YB1RncRtS+WnrB8Qk1ZStEaxEK0kZBfr8
dw6hnOSq/6pLxZ8IxAOj4hvLvWRGshkd7Uu/OAD+dpfLgTtAzqsl/7etcameWR0R
5N8X61JEgQMZtRF5gNQT8J4fAtDFNnsL2F/rsPi76R7tw6uDcBQQbg7RAOSovE7C
qIV32uDV899SbkfM2nVyCteeb74lxG1pOec2TrHncYvxN4iJZtL/Rf3io7I1Ekmj
fX4UP7eAhPmOYtmens6EJrxRoCv15pnVa6R6Kwl0bnt5Pur96ptu3JtWqlhWDX9n
kRtwYV37+ojABgyqZBXX4JDYC5oNPZ9QuqLGjqViz18ZAYTIxoX8+pGsXxpvU9Y4
f8VxdlVnrt6ATsID6nsxYh1MdKmavRyIgGOXE2u9ZPaqNF7YoxaqA1dyXXWdXtcP
+f4n8lfm/No3Ejn42dltci4xGQdC7J9JkX6WJrvjtPhvz6Jwc9jZISRH0MNVMVPX
wIoXwwNfmGgnnJA6s6A4AZjnelU46Oy6dyTQSP/0a1QM+pXMSZEgFUenbQWj7hqX
Wvatsqs27TDy38l1ywYcpAmq+eKH5+RnXBurPQMVIW3sHzcnfEQph65NYYX5hbIH
raDT5v7ZRyNpMiXTUAsA2CyVtEjEJEtm5YZNf55o96pPmVU8HuAGzk44Q7HSvvjK
vyXApoT1W4N1RuBYU9U8dhqagKCdbE8xoYAWMp4FoO7MIzGYZ1DILjae+mOXrnss
JeuN97p6KKUzLcGcgzLDIk1iAFoc72cqvFK9drZoQo0XwJKx38Wcaqn37rz7Lexy
SRv/anUuOHDqUcq8dIGcPQhwxwJXxqJ91EA8NXVYsDiPvpJVWOcomFv2pk7dNZcg
hg3WuXLmuRZepgntej11p6+7AMbdudm2sCTavs4dJ0BMUsxaNx3S5N/67RxE9oMC
CIDCjZo7kDLeZEtwyg9cYCTyzfbVavQQUIDIgT+mvQT7wr/QWOB1ftQvOuXiVa67
QA13YU6CkuAWlJRYnh+6qzPibt3VR6lAqcOMi1WKVJSV2B+4crz56CT5Zwq5vYoU
wuL1bXPtnFfMkSKrggVQl/+cN1ZgEQ3in74CJ3Vw3HsvB7pd1T73zzv3VXcOdI3O
u3SSizMBQMusgOVUHWr2i4y0IbTr+oRQO2T5gBH+51KA5hNFnh65eQKb3hQoPYW3
B/N+PBmGA5+SJlToL/KF7t3YZ6Vu6LsjJjPKGhYMlIRYCkQw2D43kmpM4OCo2lly
iPp2op3NnOeFWzM4Xyu688RoGI7OB+Zg2eezYWm7Hh1iWHyOcnt53AYqFqnpBSQS
zDTJ6XuoCPXLZJP7Pd3Gj1kSF8eHcVFZA7AlxCWZhshTVIGKPlTXdM584sWp/wdz
ATnmL9neC0M15GsxXQAIFKMNQaguiBbWneh8DyXGXqfYk6kGZvZAbRVHkh77zk3u
VUteBZobJ3MprTDGsuPSHPXFAO8qhoD804KwHBxRrKtMW7Zoy3kudx/FRbauLd7r
APHF+b5vGRYpXSqu2tjyxXwg/XvtrxURfhO+FO5H882avafMr1+Z/qvsPqHSERUK
f3VMQQSukTXJbM44L+q5LoaGjeRnIJxbszynqd/tlm4j3CJ5WRukHX0IPtkg0pLC
IG8D4Apf/9bjLo53NfadUu058eaBMWOBU/fHPtq0qCpZIvVeLe2AZs9Ew2FMZS4l
ftv+fhJqhwaCGJVqpS1hTQ1V3cmWfQhCQtsBZmQCEWihmt04QGy/hrXfSDSWUbTA
/baowsUYXYuvBIsCkhb5JyEhycPPBcEiU5eSSZFglJITOxHtkJolm+s+2TEtQIs5
+S5A0MhBqLT3dUCc7fObRDt+r8y/mzn++ezgc4DYT9MzbepTYKuj+xZJUbhzA7OA
JSOttkM54OGnXMqM1j+WKWQyW3MwEp3JNjWU4BMvefH+TdWpUADDNppjyPCNMDLJ
+r5fBoD6WKN1rXsDfA36zVAbqkMmLk9V0B+5ia8L2kbmp5TDEo4rD/zhpjvTD7Cm
ExjsPFhM/pMOo2kvG8xgLmqBUuOWrVTdjF2VppN83okgdDwVGbxxv7v49iwMxS6S
GyBlokp+0fhlpOVC2CwokCWUpugZudlF5i5lJh5sSrz7EgsT9QswSEBrwkNw99y/
/2A9c2F0XSztHgYrASvhNffZtyG7JM49Nt86zesQNq2NeZM7ggzW5WLfoU2S9+WN
6r6fPArR4vm4eg+hMuT9Z0kJmsWUPxBRVpk10InlUIH08hl+X3m9xzPO3JnqALoC
0YvaGGx8GcrAYIfMAYvMW3OCCVSzZv3gl0XMW1QFhMhIfrdW0x2KUh88GOEh5GHK
pYN+uomQllu2qcWKrIkfbP9A3w10FTeDZSeyEVpmyP33UEEWDhElbFRwhDJk9cfO
VKDLrAldf3PXmqOnME+URHZqaqKlizz+vtEZQBLeMj0qzHOMBKfxLyVvxggjzbP0
u9mQqFdigeeKxsifoYI5rOjf9i9olE7KJrxCsQCwuEP2CIoMNz9AFrBzv/Djx0Na
ijc5wQ77pFaI1gim8SnJi7HKL3oj3gQNfuKzf3wxDWVjdHJhF76a8N3V/JB1730G
GIl9oOnKqEvSfMYAdnUSaFvsVRlo1gK1Ext3VWPguZ9WGetQwTAqFpMmZ/bPvwhn
XLHR6Z2V3y+0f/IJ8ZHs82RjjqaCE2JBgIySDEAIPufW7hvgkxE5JjZxi/XxYFq0
+giCFLxwZ/2UmI/GFsxK44L12ootki9KlUGZE5IPyF6HovSlXSvayJFz60KRfFxk
s/5y30hxxN+ikSx2udU0sGCAPqVCiBdFH+6CpeqASYBe55WbGuSsa5dRep20qXKo
1Butoat0W0hfRji5JGUtSwD/v1IWJ34gNWigkIhmzpoMTw0UFro7Q9q5MXMQCpfQ
HzRAjQ6tvJ2MEODTSvXdhTRaKCK7/2AB4xwvckNc2eShU3Yfvh9AN4Qx6XSoJr8u
O0cOPsnRtTsQ7zHd24ksAzSGP0i1cawwfpgsocphGCmbockU5n+QEMnJ4q+6RHQJ
JUuy1tRGDU4YizpsJ8SFpbC6Fo2ZNG/pGbuQHH1R8dKXqx7fT+0vOol6LoCOk16G
D9tiUlF5F+OPvblzvE85F7yuwyYenfUiViMshvEUx0mfaVVLSWGljVSCsPTg+yGn
uACUdoxm9JQw1JBvwdb50aoDu5SfnZUzTmmJ0OQuppbYaLvgZZl8Gu0Q7/8WKr6n
9ZPVThikC2AVjCOueRqpS0hLg5m7wAlw4nJKcqbC4Wm1mU1gwxwd6sC9vWtD6MIw
a/mpnXx6gLv9YnuEeWXmhRNossVxextpGXBIad/6XGlbEx412IKguGfuSohuKXqW
04wbdcQr9JThT6wELZ5DX38h3M/pd2tGrhRe/MME5/8y3kTCSuoBllfFkGGgspYC
c0YLevwB5vPBphnA5c/sflBOpLiWHOGQxrUMxWDIyvAjn8EO3ZXS6o4JmD8nF0Fg
lJ8kbmONgGsadPh3rb6sF8vU4MVozGIRIpOAA5GZa2dUQc0riDneC/VRR+Hph4L4
yFAE7e7g0lEo4+A63VtDbPRvtEat2stdhVwYev+n7koJ8LoeIYwxX6GOcWg+QFcS
D96dJLUwgt9bfgZ7qpj77eKUERsgZe8NKEYpRVNi+U1IvVghPtVjNAtk/EwOxCrk
H4n5afli2x3aQHa2I6USq2Vp6MfdDsH0hF52Lj72r7RpCQYg2esmntQWahDL6Zzz
VHjFGw7TvMlf6AEEn6QGvpsBwG4Sn/zv2Qm2brlFOI6VV86IRBLj1x3HHdG1LTJe
nZpG++L2Rzy3zJDBtvct3/uShq1DgCyLKT6ruDkgto5ydwzQvI380tz/RNxf2nxz
GaUqPz40sPZsBxIZjvQHbU938/FjGTMLypTvL8ZgJBNhPWNXkRw+N6T5cdjXvfna
XqE/PlkPbfm4sZ9r1Mredv+1YLVilm+MYvhxgFcFyibG6M4rT4Izex1eYDiU+XmW
ODP+9kSO4R4YlN3C4W5WAdGqqmV0nf0H7mL0DDjna2+oxy2qCNYNn8kS/hvl1CZq
r1NZ/bexKZ+ReoasYuH9cBzBEKMcUae1G+ZyP/3AZQpGYCop9MyZjczX+RtrALER
olhBhWHma3uujzk6b/2YJGQk3w2c+bwV80CzuSr+GGf8CxnrMMHbBvWWFVGmio92
JNfLi6DdyFZLW29hBbvBSweptd3eyMLTVrH6SM/gxflCkpAbRybTN9X3AYlhIwWM
wC3X+bnQUAVZKjGNA+aTVoIPy6bY3+6taUrftxxjqlevNXArmyNXu784gd45V2rw
mIvp0RloZZCwHFr/higxdUcxHgrSs8/iu7unKkxYb8zPbFJEV3ueQdeL+fik5qCz
8EC5YL0v/KnTzio3Man4TGaym9lrbAXnb2UjLPE6eX/LjTydwcpwBfNBPlCd+mTp
wVDbWtDOcrAQ8g9sJso9edZ4d+R0XGgD26GMgoM7FTIW9lM1xENkZbrO//Iy2rSk
o29cofZds3l2t1SktUcwsdCc18JzmlEtZNfKeTCtRrMWOmsnRGsXBH3T+fWt+JRw
r3VheIyYN4dE8EiWYNtiTUDHkQJt1jLu8550EiJonwitPsgOOrlUZf3ETOk0Kv/g
TbDqtxDWVEhZWtr93Ld9A36BfRRAEQ20wnM+VViN+KBcpEYAL4BVVBKvU8KTqTDx
Kxu3OIDdgorwkt/2Sc5AbRBf1VMwBNQDi74woD74XCyViNOzsNMwKgyXhXfQAEta
0ZipMtvzSbl9GdlPlObmo7FIJ4lXQiuu1InJL7Au23VPFOg69VpKBFjFP4IC/QpV
cZrpPbp1ptMi49+8O3QCEWB2FoJvRGb1E3aUP26GPcbxbUspWrMULWb4TNcphnSp
qCZt/A0Do/hef95Ze3yh01HDxU3nQmAvGWmNmHj+R2q6u67sDD25jhD72+VxxO/8
hoO6Av4C7dPj2TrNRvz8+c0KtXYUj6DpxsoRU67TR2tvMi42pMrjHnlf6NJOF7iU
tsn1CfUacogcmyuVM24PcxULjAzzDxgi+iNAT9WCsUGroxEF+ZdinCo/60xYhFzZ
nheDVUX3GKKegKMio11V1E7xNf7OQRr5dnqRWq3bGmz7qcHX129SFCwgkRtSSrmw
BFG/QAjP/WUTVP3u+9/lsWXny2iNTMAuSjvnFZ0vCy7kclIq4I8NcyMZZHQ5XmUp
3z0AWepE93smB298fzXs9W42ayjsoBhE2tyytzLeSCERomy/iB7DhEtK54RLDulV
y4a3BICUTPPrkefAv89g3JX3Lt0QbSYRA04sk5eC3pA+jeIAYRlKK7SkxwktUJR+
/Zv7rsYdtnl4UzTxmhZdrryJWAFxa3jM8ogUO54mjhqrKxotFee1nO08ZBcPFdtE
7ZvPBYnINClzeSlo1x1hzvD+/6lU5PHCkt1WZ2SFmCDbhlfSF03obnhD7epKc1n0
IANUfcs+wyFID5fwxPnn2fDogkYJ0PP+onbg60asTmqwmWw0s14P3vHi+hPsx0gX
cDiw4MhENHHVjfOSra6w4Qj2vHbiFcT//34YnV14utH7FksVlhbDIqK/a5B86Dqi
M5Wnc/MCasHliynD29WIbA4V+I/DbHqgTeY4/amGzeemidrerQDNwEUc0k2ZXA8Q
D9rdTV+r8x8V8NwFxeEpoiyG8J/iFhLwnDOuoKLyVDbRnLDrd/fOhZvrz0QqkKiv
26K+X3ELRZaOjn7LFOhg6tGSm5MqAfMrrEn1I3e5GCE40vERaHXnO8CtBAQdjNst
W2wT82OfGUIlwHAtNzddIpPryYynzVmbg8Qz4X26V6F1jydsR7IrsCfCeuC9b9eP
Sx88m8dnWuiClIQtitdCMDFAS/WSmk/ePJyMv9kObGqTxoBHnK/B+iyKsk2klqvF
0pLFY3AcELEjxz/es117V7AIvyQ6avTnK3yzRaLLumbWVI+t1lkB1ri2tF5Q2Hw0
tPdu6nkqOqjProzctsjkb2xX/qI1obA+SMKNxJqErLCM0tmsURpSik+DCaEoMEib
/owZsCancNXozrEoyxGXNou6BcT2ujhvFzTuDplAB1rn7Omj/xGUeu7mVctgp3AT
JCJwydrOtzIjQf+CYRHhugkGyC0RZSQHXgwvjnIi6EXpTfkAysFwxDBqpLlW0uEH
kip1HY9QMD3OzuFgof8FdoX047BN1i0CvjPMrQxZhZkv2wHjgWnveouJi3olf8Fb
mIl40yEie6O6QdvVrfwLFGp3nv6t4k/JSK5aMn6/euUuhOAf4byJzLmPruDBtoUA
1yTEV7U/XPkLAWeFZ5FQc9ZNkIvYtOMZDz5o74766OCVZi8ob0sCDvjpm66zk5fH
YIAORCunf8B8eoGGjvaKWeofpQJC9EQTw2N+qNu+tya053uCnRQ+mL35ObXvYxd5
PTMOG3VSypPjy+Msdi+CutSRPxwFrSigoxnkLNAMVEyrxXIMvdY1UBmgDIgp+hDi
wqfLNtK7pWLBb1jIc8LVcoE4CTNLDi7iMqYa/5ALJfkRqY3escp1at22bivvftah
FmmqpPzyHOCUFUoha+apG6gLDacOuaBsaD7UBhRN2wk+W5KpJ6Iod+iYiZY1GWGF
oj+7M4TUYQlUcM6Lp1GA6h6LNstTr0RFddc8kAqJQbzA5efbr5uyyfjK9r5GPTAl
0fCNVxumCRkOI76KEtkPrF2ilwc96ALKpzLQY+A7eU3AFINpQ1LzZukVB4CyjrBv
qWi4wSNRzrvl6wLCMYd/Ng1VRpUhwKz7eBlzjeYmV/gSRZEh0RCFySdqjdlsYc/1
JRh93TT+Z2OItDnNnuWr67rSZS1gYdn39JohLBRgMz20Z/fsz2HIYJH490XQ0xym
swhnSao1NjEYnYgTMhHXruyiUGxqjXknfvg3/oWcne8ScK2Jva3pHP4HbRlFMAxt
F3vkhXOkPTum7Mw/Id5X+6Gc27FehlfhVODqik3PqtZeKC1ulVu6q5C9XrtPV18g
hvWcOjMkYYRgN97RUYQkpJFooFA5NjeiJXgFAyKRD/ml253McKo79m1tG7BhbbQ1
2R+RIfwu4BtV0aIpQKPgG0A9l/PI2MtLIc9DBCnN/qi345d206BgVzYu29g1J/BG
WzqehnBknecnpz28ZwHASg304xMhi4NbXiFyjEsW49S8yc3otrezxfQ+y5CBx5aL
Uyt99RdNrBgbipZnDCF8qr4LcM1eirP+f20K0BRYNZ0F+VznmWqoe152Zp4lDPXN
ljSQ+Qqf561I7mAciBTMVKzC3c1FQYdzKGP7L8Yn4lRl1JgiL1tTPySTxQBTaZ4Y
pIYYqFPDUpOnFHR89wAnt1srchlEG2X2Xs1sFlne2+/wZFDOaAI8Um3Juvx33LAR
ib4F2qcKxnDdf5+JaF02AfQnxTIbgwxDLMw2EpYSh5UPdd2u+/f2BneOj69eAeW6
BcNP2JFESn4oKq5g5tyV+wYFQ9PRV7wPd19mzoNyBdAar43Pw15Y8osuT3iaUw40
iKLDuSt9GujSagFNicjInpy4VLeJhp4V3L0uOdd7wOmJGcXGETsYbqN8H9A1kYcw
ACalHsffr+rY3yJdWXtC4F7qbEmvE50ER6zl79uA3PDCZDqqCpZ0onk8DXFqkl5C
Ogb9TvTaBgqw6iB0Tjq6qaukrrxHSKSS0bEuivql+K9BMGA/G+uzEmTe+MNLA5Im
vHZk1Tk6JwVRNBTtrviRVKwXGIka/rElBAy7NLNZZ1wmoX8yHwbFYbEWMRZ11TUU
QZmW9AixXaa/GTY1kbUKNals89gPPuYH2Z5L9VrY6O52MMiuLnW3/YB7C/sIuBPh
KtsKJslJq7mTV9uY6gtV3kT1VW+5HVMHt6PNVL46D5ZiD1qnR/5mXvfDRC7/opYL
qGv24q3MTjwIZthDLHF6WQYYwE6Hv7UoPcGPgXcAdzmgtyXMK+teOC0/X5MKzxjw
i5Kp1WFqrz96y74rR0k/R6B2nwjpw4oBKgwaulkZa8tQAMypABGXr9uawPmTjuul
3S6jFNQ3e7169KyRhAIe6C8Z0+J347PS8kFWsJrFNNqIfmN3y6CbbfN1Re3pYRr8
NSuI1UqRtVzMP4NGFpGpNwwgSEO+lUTxb8e7ANTzc1X0IvfVUhpxCOmcFyF7ddG8
wamKpYZv5NCt7/dSBcAvScbCc5bEf0Upbn57Zw8l+XHSWfT8M2Y/XjkaStP0rMgW
5KmLSKqUU3k5WXhOo8MDsZ1rG48Vo4A47pY/skMnX3VWEYtg0vTThkf1erz1X7Wn
F0evAiKqohxB8fEee9QELSSPH21dtRsf9wMY1nilBJK7tEe3StzAsK1HsKoyJbx6
sDrMlYcTCs87fcMBy2qV2HE7Cl5LnMNXohqJP8I5qx/SjeCOZ4NnuVIPLA5J4Za8
a6wX3qfk3MW7l+l6GOhYAWmZJXEwGkuW+rOkpNfV36b8DD/O6+uhmEYnAlaLEy4Y
Fd+PRnmfKpkT1Ko6D3ohpMnL71gdQ8TXdgUQwj78rf+LHbfCwnHArq7QtFFBuVp0
w5H2zCdZQw58qwl3eyKXEta5Po7hxVHmiBSk65Wj5dcQ51P780oYbPuCYwbxmBmq
L/EUh3Yej0IfmvZmUK1KV3KbwBSVLHM20pxJU8425ujLSnUT4X0dtkWj8HkhPUuU
jtj9xIPXGR77/Urff+fG9f++Cgi0v3+04XrULc83euUUTTNX+MgOf9M/D1xadUg4
yvvOkdRugD37aYn/fZFsxQCBMwaehUJQzR2bk5WMnNEU8uK2NBct/UYr7eFD/y7d
+hdpf8jfPYcqRVZWHF7CTXg90Fz3+23/iyuaR8nbp0JslSGQyVO9m20V48kmBBAD
WsR5BuMsIfEPHDxQ2EAJfO/qHQbORAl1RltcsEk3tBZ8OP346E7+ArppSevHcolw
M3NpmX7VfrojlGk3Vy2wYciDtMfeS+gwa57vcJQnCp5Qr9MtVPxFizzyAfUNfWQf
zdqTelqj4l6Ls3SHgqgVKEr1XdbA5uMeGOu3YuYxhiPH/SgP367Ka73nmSy8awDA
XbU1HK7NtJZom8C96HMzuFkqkkQ3Bc/Un5ZZD7JZ1oRqN5mrAKctDHZe6yjcFqt1
rVXdnH+QIcSlcDwqkD8IkhVUqCS3ZWZ24NHWahcXEhBOtHY6KfGr6DbgP3FywDjb
3ZaKUEdIPBlaq++DPUGuoEsTOMSiSzQ1Dq9uGdM1L6xchxhdO1DuyLzSsfl8NatU
Hbb+j3/XnetOzrEEzIRcyGv9iIu3a6qrRzxPdrpcvcS/T6VzWhKFfYQhr2QAHVaw
6Ae5mn9EzMMu7XB+2UYeThdCGV+N5J/wHxSdn8TPydJDDpqroQuHlTwl+jLc5c5s
GE8+sasSAZoV/0JJDDhhXFRxWBy5FElgQPBuZejrHnqEfXXnccXcN6m6zcW8FRgh
jUKceGVk18ImhN9E2+l+qhrbgs2XMBLzKRdGFN7TBfZspEP7tumKd8tcIxq2ei1n
QmQJIcXWNl/NyENUwoQz1DhRtnsK8Y03KRbsn/+N0yYXn45Ftr65p1/G3UwZ8Cfc
nBBdb1KpAoBK04gqDxzCLcZqLvtG01CTj7n94lA/OWzdal72nfPP1BupxVIzSbdj
/bGb+Bfgt95NV4lelUggCztpb+Qz183SdtftY1TEYDGPqFWYbHe6OSQUD8uHYt5v
tZAlQALb2yPH3uGsf8skwpfHvBt9O/OEwLRVFHE+GkrW9NfU78Q0x2Xz2RKN310H
dFZv89omj/7noFss2gMiz/MHU29BrZSQD070jJ0uCh2vosokB+0jGIgFijw/awzR
ppvyA/gcCdp5QXm99OgDg0PNC2bKBXQSvh/W0Zw2nnWFAqVigcVeOC/ksRFuJCId
v7WS5yd8hrrQ5+kIUqKXiicgzmUNAK+CbYf1X/5XYN20dQfHGPBOddgxh9gNrXs+
UcurxSMmNFMB7also3ofo06Tw9NGhjEAoPCuX8ealyitwcjVYnJDuxx7mNokT81q
Lt6E51px6r1C+x9mRYiRZSmIpldsY75MZI5NkKAjALzDm/tHg5y1kxD70SaLV/JW
sZcWWc/jDyWPLDqPaycae4jFhPX9DHcDV9zkV9OZx1/YTbzQo6lwMYgTd3UMS/M2
Uercq4DYC1MKDCablua4gUDczMxydT4CyIDOFx0HJuvUz6ta4t2nNOeR8FtcNFiq
HZLzkoP7NwYOFaOKDDDOFDlZDKqXszvbTMYWLf3FVD+kLAFTeH+6ajasVH/ZGqgV
R/VKCVmdcBOMpxQionU1d63octLov2vC9FFYtmSmFDvTRyTLkh2LJ5doesHUhRWN
U4xIqWnZtSIqlj1Ck8JQy7F/B6Zy6Qs0csJFa2iAyx0ar0HfhTF0e0IBy9M7JLfP
VrOdvzZ0TUacuInQflhvn3IpQ70ay92J2WrBGNmA1FoD3Z1YgTdsCnaCKiupiP7K
qsHRoCRmLGDE2Rqi0ryKPr/1lwG/KOIp+/COBXz4MGSJ5jBw0x4fnnEysi5242mk
2suVtOagsgHOCN3Q0QE/rxk6BBxE8rnp5J+kUfI8AVFDmSoB6CI/eCABnmcy/o4w
jFLUYNgPNwura3n9ZAeK+pZMReS8hxph80Kzjw3W7OD9EOlKBBNLAptZs2x/wY0B
9JoOo0H/iPRWP3llR4Yi4hL/kwU5jBvKsI11Zj1Ng8PyV3m5VxFdaUhux8EkWEWM
xL1inwtqQMzwc3BCHtHb4unJckqWXblDPEgjJdYEBqBrJGH/uyieKQjL8tkzKGX1
yWvXKEs/9VOwEXi00G+c5fF9pG69fqxIH3kpvRtTPGl0rStAkqVilQKxwxmbUsGU
s/qNxGijX8RUTw7MTVBeNifLiZJZQVpnI8cjdvavreWgs6H3QEkaksUj+zXZ6mqA
7Emi4H8yCvcLbLNgpY5qyX5iQerz0vamXph2snNervpkMCvACpgXsrbeYizZctqQ
xBiCZMBZIkmwAXbf11z5e9M7nI7jh3nEJWB+AsWlrK04sq7feevxpHdLPw718knA
kwukto8dTcHJjOkBzyx/TgIGbrTlUzUfuJWXDi/fBGSv3qDUVY6zjHMsNYprdtSG
mG2QM7Jn+NdKoPSmzp35gLamEh6XuXo/4pFbbUZQPpY69thMmfHiy1BekIvCVXxd
obelYF6tkXpu/cGx9NzzZw/ZyEEBI5Ghs+Qw1OFBsZvw4T1b3wE3YoczE0FD8wiE
jpXQOQsY09AXX4ASDjcEqSOch6KNUJPZiuB/HGzETMoyj0LldIqTBXrlZhLGTzwF
LK2O5Fz0ZdnAk4i2pYn+7YEkMwPp5/qsk7MrBQyCrcCKGdKKlcRC6McxKYXpQyS8
QEn8Md10Dktd8jrLnwlVIk5xUlL0VsMVRedrwzGlTYZzMDH4q1m8PPHCrRrWvYhi
gNfuTEu9oEbLxu5kXr9v+Q8Pb8WC0eJXcowv0UPC5VTa4E6lx+pgDWjfWCrpy4Nm
jslopM50ocOVEhFyP+/TCxfe9q4/4ShFuPHpj/Y1tmxk9hkK+sGWE2cD+Wcyk183
0CQ/RSn/SI9mbY5wDY/VHCUEfX9fex6TVgTegIdKgdqVWPZxnyjgGDLNrce6JEDj
7pKm6peQIJfjmPdGeWA79iA6po3SX81qBWRdaHUpzBA4SrF6aTCCKqodqdewJKy1
31N63flFkI/fsMyb+Hh5I91zL+ChrD+yqZha6/HhipfIyOwIGApJ6gE3sTrR49j1
S5bJ9WvWcZmlOGfviMOZ9KIhFNC778Fi7veREK7lb+3ppMIH71Op41MPDN0vP8Ah
wUgG/B/252njIjUYvM9fUWUR4jAt4DKepwUhyfCEpPUpvLgOabfbjKqS/PD2so12
9y1/2UBkRMGJ7uuPyig9gwhpO6irrJ28HSndvY9hFax4JbKBbatB0I6K4Jg4Wgid
2yz5Vadnwf8yldNxld2rkVzn1sgy//UXUZiwVFW3Dt7UzAAbHrJMwW93zmeuo01h
KIdfUd1aPYCBzd0RrcNqnCsZGZzRrQzWVYir9huqn8ffctmv0Zo3h3j6BjOq5h+f
De0hfy5IPrMl5kT1K1za2RQh5+u6ogttz3NjttlzFavNvXq29O3z5hZvbuFyrvMD
xC6U7G561Rx5eeszpjxwlaMrfoLqxWK+EjYWISMMJxd9v31cydv6OBpq02IESysd
52gutso/vLjBh+srBWvLt1gYTrN/t0qt/bJ30C9aHmGI4OXCG+EMkxK/bp9wXqzV
ktyyXBatuAvjYPURL83IvawFw3BNIFQEbV7yeoFu4FaC4pABpv5UkA4COTKrR3IY
Z+lqvHhCLwIBjTzuTcw7qyszPjeuRUtbX6MnCu0Ga4VRUe0dRkLwQjkCMRetxNN8
j7hQG4vJSdgW/p3W89VmDWPwQlNBEqCCLQac44qOCMC1NcFhEA01JqeWfhnkLtj6
Gy5A3Mu613taS3UgQh1AIHav+IiveKJ7+JUf+KSRdCCtjmd7T3CGFSTy3+WzC0M6
y6A5yX53T7nyK7gLDJJoAXRmZv+hD6BoKxn8mKgHVhaFMs9NId/HncM8n809m42A
CS1ZvsReSpOipsFj8VEA/9W+kvElLwe/U5YF4jG18ADyuefpJvr/ub3n3oQnN0o2
JT0L9CDrrvcpAQbvAY73AFBnnkg7zMPJK5+eXCRnn1cOqn1AY7knG5lkulyNcrLY
oHEOX86BaUwmamsHqZMF4PNZaY8ktsmG3kcSH+KWmjLhLeqDPoWg5Q48/aSXmEs6
3DbytQS5hLLjqHoCzgsPCnPm7ac4u/E7oWjiWKBq8SN8CxzddslBU66gaN1MhPrD
qtXQaP3Nli8g1+leUwYwcw81q1ENl2q/HZJugxCkWwXGQXpDuWZeEGfgCyMlu+St
RcFFCOxk0ULwsXzrGnE/fj7IuLi2LynaP2fTsBlwTMZKeGEtroT7538tDES4vPMS
RFmHhyR+MXkHya8vgGstHvwHnhHk0dNJ3E7eUlfBcH7gU7G/zVcnWXwpKhr0qnpH
Dr2lglecxcwnWZBiAp9B7NaIxKbFbmdzaSsTaNH5YhiJ5/tY9XhmUX5cVHHECKyL
nSoSW+gFal+G7cnq8gtkgy1B/PzUafEtejJPAjhNPc6TEtwZthHCjYc2HVLQwyoT
UqIypVLBvmYc4Aau4QFTwE5DKXndPfFwTXbDesNiWSAbYTzKpW8NFPevPWZt8nG4
m7482Q3yqVIRfuYJiF+8jdcjcP92MQzcJdlUYb5s99qD3QiElua/3ahTX5UddoQm
PzfpAVWL4JSILp8loHdSOxU3qEgsAiROqBM/DKHasasmrWRAhZzee7pfIdYsTM4C
+Y7Zna243F9XrBn8ZKvOz7yiLR9UdxdZr5O4R0dOPkgPHFp33pNHlUgpIScZLmL+
jeFaLjf7ZKYptfHCgT3QrDos8pxNzdBBPoLnaG8sfmlWskm5FqT8wsmxqaBVSX0M
tiWAcWYPgl/kUrLoU602AazCyF+AWrhoghgbRv9sDVslQ1vJQWsrYVbBfu1m9TsR
H8+9pSmLTmFfFOBVf5P65a0ZGq9vm3nN0tiNJ5gwx8UwIHdpM5FPKbno4QlVSLM6
HhzH9y6OkFVIiBXskzE5wS76OdiCC5CGEDa+qjXSjJzXZMPCmiP1BZfwOljIaw5B
wbEvp9VhRDK8J4R5Qmws3xBVhNK4PlTF2tWarvtrtFzegjEp13YBSw7wBuxlCbce
dI6v2Y8+kax/cLfZtCy1GLrC2xjPbM+Tv+vuCpyPwSqVo6ZOpG35k2mtyvMFLbHk
0gLt609wJjUpSSM554u7VSM81Lcc0K+pTlVeHIqT3Ov09QVa1x56sSAYSbLtHYkB
vLE4CsMGtDSeHYl5GhgFnPA4cAeY83jb1o0bbWq3zsUWddcK5d2kf36zZxUKZM+M
qjysRcGIH3v0nVACYe1TOi8NEz8ktZxQQA/oW7r5OwybBAYIbtu70CFtC90xxdxL
PLFUJOs/kDIh3usI69erw2X4TiaiSmVEoAh03YEqxqTA580H9XqjtTsTgI6WmOL9
HfmuNbXLxrbSBnld9D8RVQWhzt90gVuoNcDlU8bd2Et61g0oqLqliGVCs56YRYcU
D1dbDfeU+EtvT6iX2ySpbN7WUYcjc0Nikq/HVIpiMZY8a33fZHXQZtPTI3+1USCV
JpEtOWt/gHWMD7QrSc1uCcuCWNpAyl0Qy/g663cpRX2x9eugX31IPktJ/W/Ai3Ww
1oDwEeBxd0JRNaihGD2Zi/cpNzZ57n7oKLGaRKHD3YPoMhOGKo87gi1/dHaIDqzB
ovWnSIvr9Hu3zvOe+vOwEnfdD/4jGSbncuA3mR9vjmfWfQ8TTf5wzemDYL/KszWJ
OUfJaP56XouAUBJQ+Zr3J9WFrns2VYbqZN3oqU/jhoOPgBCu7f5MypqkkEDjv43u
I4w9RlxUKFpOYFLHXB9i6bZDZnoaEYF7A1wZgt4cKmB3MfSLp1UkaFgcu4ny2oG+
aqlgU6IZmQVwHTFRyezD/Y8Z/4GhjB5EAjF41E7L94w5sevMJOoxoiNSm9PeznVr
xN6LC4csOJBcSuE3bEmlEcGzVdqlW0oXwwyWWoYdkXKB5OsIe1c2q8EiA0nAFe+Y
KcCVAqXC2PONKLsgRK+o4v3AWzd2VNgKB5ExguHl3JhNa58XQxhP6AiQJCwk8biG
RlSqHu/nZI5OgLtFYso+D4mkp3nooBxrqhCceODoxv4pCt/l9PcXQEmuDA4tLnyW
to8sacUKjM9hnEivmEmrk7aQig+LVsAqVLnCBBbyejfNVqp+13uTRMVKrW8IbgAp
4Iw2juQt+XQ8Z+Tit86cAChFEKkjR6csI2diCV7v/oAHiMxGG1FkFl36XXBAjXJM
ptt0FbBqNtcJDR4rRHyVGlgV/G6kE230sMAvlFpG0enwszoTw+oZ0DGsU3RWHAj3
+ISKazr8aZRiieG0/4sjpg3x2eAifmPozKkWzZSGo9FHa7ldlJrgmJIp02YnRbB0
mAGQoORy865N8Al3yNB5xMwYvdGhZ8j0ZlpWA+vwS1ZPbNUe4vMR3NP+tnD5gRFC
l1/laU/NnWlx15TFQmh/xGXN0DQIxh8aoMYe7o5uvubEQmFWqbJrLnmPoajdx4pD
1AvlYC+x2KDtPcyG02VzIroTB5fQFVPUfXdoftREPjIvLLdPaNsinlPJTW7TZHvk
4uZ+agoMB8aTNJ8pBNtXX5XvvI7GafHaWFzFkODiR3PzU0GveDPpAGgSQUAzKReK
+lXPq7QF+RJNHZ2qSzNPXpUVHj/Uo1COV4p7ZtMyQd0WMm54ZRzC2hhd680Hi8Ih
AbSzUqYU0Nd6O9ZogGe6ru/jTqYddGYwWBX4Sm74ZI7yhLn5YXfnj1TdzLmIWeX/
4keiQgEcUR+lMp/F3nvLodLHy9MDp47UTfMomZ3ISOQaX8zb4F6VAsJh4IB6zpCg
xEgxFfYKf6fiZ2pxcUjlPi4AufthLyNx+Tvm2/lqfDtOgtXf8o1GsN+ZYhq/Iof4
nCY3aO6oC9VXSk5XQ4Q872e+zd7F2ukX+QxylKBsdH8DU224K7LhqS9jVA6tvtiX
YxypaI90yBN83LgQwkiRT00H7LQ2lYL49wXrTkybmOXE+ULhH42eQxIhmW+lXByS
ZYPoZJ5QJd+zyQHyr1LtYYP9HOHFkzrfNiXu7oXt2TYJseDNPt3fgry7UInm3s90
ef37v4TOCCF3pohzhEGJn9uUm/TBBoo00JoiUO66to808sNXiM4oU9VKq+ZS7cGd
J1wwJW1u9kPHtqrnV4mIAc3m3DkGU0Y1fsZAotmewiXBCzbs1ptL/6ebXokYIWHc
9rhhOcZI/FQu4z7eaaq9G15B2xPSdR0MSlqmzGfSOJbduy4kPsr5QhQRvcrge18T
WxKM2vzaunQqqdIrC+vUh5G9B290r+/4QgcVBPsC6mRevf0mbl08shat8gErzZuU
1Pfqd9YXV0/tcysbPWlNeqXsQ1LNOw5lwEKpNUB69Y6UuajPsYl0YXN7IcqoAC0Z
KwdH/wXVlsxjQvHqtz8Ctay6TI3peJqxf/6gB8bBuyX6jBcLE/0Gx969DRsKEpJ6
H02tORcvlmtvdzFRZ4e3T6cKOevenzWWGLLteMd2n0A9Y8r1j1JCvrgYXGEUtBHf
xTyEW4Kg7mjUzCfwnasb3GgdUioxGIChDWb12OWwXMXZoMppoHPgKPrYTXLGny2E
R3x9ZjyLOaVGFmgof5GzygVKuOAmyRnNED99dsnqkCeuoyMQJAG4thShtbMxky1H
8sh4dOCNegC1O98jm4K5InHPoNIeJfv9P91kekH0Bw2gkdGdwqB26ucu5T19JrTK
VfJBL+4Il3Lnw45sfuvKAlz6vTEfaKy9bT1dVC1dw+9PwqSnIN98F+tU3qbpnNNu
o8zJt6gOVBw1rG1rt6USAT56NSNIijxSU+ovv2VhgsBJGxW8co1juXsruMNv7u/W
Ct+AI4OyzEMk7WNY8+JWzINxmV8m7HQN+9cJMMYKo6OXzXlcTfWf+DDHux3tadZC
s33V0GA/txuhARxjTvpJ6uMPp/8GTUNdnnRWl/hyLETKjWb8xBwvy9oBr63cMkKL
7CeyqFF+SW/6KKExRnSqmSi4bSm3Mqd7yh0+gEjHNwKGAFX6CmHCmvxWwJhKxiAT
cPz+Xpw+slvE91GDqL4Cpv0IERq2n94N1Rkx5zG0ogHomKfK61gP/g06F2A5Oplz
YxEZBZCctSXWXdM6ipyyFvMlT2d981OLrbneI1ICA+nxeQ4exlJ8p1mBFT2nj9Pt
A0R6M5pBAymOi03O/kMEPCBI06SwKtLI+13w9q/m/SCLHqnqaCn+J2K1CTAICQ4n
u172U4kJJx0FwIC82qRnfynmG6qMFeZK/2UO1PHeYnONhZJvnwhZuzrHf4jmmfg1
naagaU+Ah8OAN99Bl58Vv2Du7cXVzrRBC06cmoG+GO5YMd6oZYBOup8fRNR9wIvL
gZF5QE0Wh7aeVjBecEih02lPb7EmXNRCmFobPIC7Kk0qV9WRa57KeFvnMlAOuKm+
9UHUbac5zBbOdWMIMXurSLL5x5fYLNQJbxurGW5yeX8z8UHVTRBbOvvu9ttqD+he
2t6ZWwGcem6tPyrnfE/itZm0YsizHz1OH1ZT5cR0YlqvAc4ZC1CC3CqqJBW1arbT
fa9o0Ue7UL24XKqkpE+QAQoA7l+iZVuUka7tpgdrCfvJoxLHQSAJcnzrp63zpPrF
shDWGmOOAFvWfRdmvRYinlwgZ1zkTVDn4Atoy5uuVPl0aQaG1pRzpYSyyF8MjjBT
gjugII+PXyqfgwsJ9hoH/ZBc5mgGJh3Az7lxj1NPOa3Jd5r3EKhJ4D+s4pUAyXsU
PYM9T7QkZR9k6mqPdFuOI/6Blnam1TvFENL9cep3iq8CrM4XKqIRSnBTh31UFYas
B7Cnw/cT3R1fkmSjnDwueI4kGjR7vUmXV+4Y6x3CYDbKceHfNcRLbivL/rSE7vsg
2vscKAs5eMqKhCeJo1lRwHyDnVp5JqyatcLSsv0qsQKZSxY2SlHBxUkOBRuyg1hf
XzSaY81ldtPbdR7KnpmQL7KWWMjfVhcpCXopzA0dvghO7uisOf9H1eERkquuhmGk
1krdHbpPbh4yrvMPcAHqK9+PE2Rugqlb1prVeBxZvGX9p/DZav7UR/1FEZMbX6pr
J7EUhYWD2GpsHBixhSKmzAoB8kWJro6RRn1qGKebqrnb9WaysKcIFhM/3QGCJsBa
NZgO2qdEGq38DEfsd/2gc0K+mOUKzPsHBazXz0N6VaEZ6jr/OQTKvtW7kqbE7cbs
sdqoe19jtcDk1XgkoKM1SB8JWqWLP5ZwcZXK4gmO1hXN2Qa+n8Da4AS6ORMVh7/t
K/sYGqQEM8bVBYXjVz81T4gH5EJ85ozLFKtaw//InsKA/c1DYb4zxqZSpfahkkEH
t2KtT5AKEFcAjc95gGWiqn4udJKgPE0VnU18KXnN4LC/C1b0oeUO0lS1PWAVTHPa
LH3MByqsE9h+ec2jA85WzUJmeHx99b6EuvDjTAHC1buWPv46uHGR+veIvRAJ7s5A
1Gb+XAutBdPHA2GD9vYm2O9CKLNHldeXvm4Lb8A/Zl3x6RJjYnOy65ND9dQqUjB2
C/CBrEwFPNAP8hwc/AnlIzkvb3bzk3ntH8ybT0AIuxO1mGcXOYnOsrfVdQO5SLXH
7oyLNM6DKwueLoEer7vAPfp0BqbdtO/S/JUeEVc0Arn5C2yXhbf55QcE7CuPBXVA
QlMUOadetNIZV6B5bCe/21O13XBIh2qJMMebJ/Uae4+vKAGlZYlezYoGNI5RxP5A
Vwpp26BHMa9oDwwR0/+ygG8lUSbIpaRDIj8BDwybhdcvXobUyk0WGM22E8f2V6ac
c3WLiHUy5yboeUiztxD7/C1zHhQ60SKBK1ABpyWRuMMVFS7Q4nRqfcUHfj9nDzZ/
qt/RoTycRxJfLoflNLGcPEHZRpltoP4ul/nDTWeQ4qgaa9Hsks+cwovCbvn1vQhB
pEAq9cI083jnmflXwJL4xjuDCU9bgbwqVU9SBnX03Lllb3pmWV7rfNAl6G9VqW3q
IBEvkkM/J6oMEKeOuTNpUjZZsEramvwU5UiNxc+2pfrR16PDaFv1NbyzK3O4OSfN
74nG+9/dMSIEckb7EoNnxMhzHZERXTWD0l2S9lmxYNsfNSjxXIcPAM66VfNYbx/F
7kU5C5WdYJLDrbS1JnUxA3QlR4a0pPS2/h50GWNJVhrLVXu9LV4xLMBBX4UprOHa
Uim9ZTvR4hbUSWEGcMVWPGRppq3MwlI9KGXN65Xne52l2uOBYLUsRwoEoGSlqT7s
WNS3NVsrjCqV/SKGGak+8toAiIUu7VOcLNeyLdEGP68agcWmY/aQGEku2UPGGNP2
OUZf+6u11DQ+57pXt1sP3cZkDW50US9xhCub7aNiUsno022W+RS03SbSSfmg9jyi
VHoHPzP0l5N6xndlhRaV6uIZxEpJIW+IprCHejLEg5svsChvnNBhdSFpnxbU8gqC
XyNVOg39tAtQEdbcnJhjInUEfa+CooHW3kuorXN6V5koE9LfmzpsRsCg7yRe0OXj
/UMISgWOnotYMzlTK+WcxLKCZ9o8D7VpXtrTS81t0W3vrKx9Ughvu0i0sNV+/a7x
lPDDoTGPG3yT7OpBH0mo97mU7nwcYxzPHkN1ZzA9DdRDz6mbi88DVE5D7ux0+H7/
x950xnfZcykS7CAre2oCMfGDMpwGKNIVI3Fx6gecYDf5hgoz0Tf9Q/2zsBOpBYNC
Iwv+7tpYcunPZSfWQOu2P0GnJ9xIuXGc2Vu+5c8oOpCsiNm/XuJB23RaEz6wto6d
Meu67Z48c3AxIRLj+1L+alWb10FM5tj6jf8wW6ruh7hpluvclmmgGCsnN2MyK1q3
S+ynsFxkDoOdB73rQ+7LtS3IKgfjQgNskGhmKxV/j44Lp3u57hFdK6EUhHc5LXNe
TOGSHwC6M2xqzwC4ITpG31IqpGP/sRGMV0xqfPrQkFTEs+uNbJVpja7vTJdI+zRM
6vBbSREDB+Msk7iBt+afXGwtIA3+krqBVhmcdI/lYge0/gA9YUHlyw2ex4IjQWc6
kLcxu19XgfZ44ADhVb2QHZXlIMvbgwdFWAM1yYJQMzCq259lPJPm2OHSsj8+/PFQ
iZ4XaZD+H8fmaO5x/ZbCWepknswW0oaKdVZyCa0VIIXae4VggOra6CQnTYQvJZ3d
57FZ2bhD9nuFyctZImtnmPkkuWMauuu3tmnrGC/JYBJtTJQfmok3P0vc2/HsGsn9
dMXkIIrN9clDsb29FalZGIu9e/nYcQS9KiE7PkvY3wjwSpZnc/jjo9Qtm9At/Uwk
m1CIV7iMCH8JknHvrUOagikAMsCK4eryo+vER3Kd/4nsF+0rUwhVRaSP2yYsrJLF
JAzb1Fc1Mi8qo6SBF522CGZJtIDDjc9ok5UDdTPyo3PeX2paApbYvLjpTjjIewb/
cnaDXOW+rTSI5qO59kTBDcIkN63RuEGi2PuZq/jN+z6sJAug2YDGKvE/TncQ0iNB
fdnq8dqp3gVRI2BXVwECPB4QmAE7Wc7NGbsgKbOoguHvsE1LsrtVg0t3gv9z2QWB
4oUVEef8cvn4Ne/h1c+y3FcD+MhmeyhoVc0S27jfKgz/xQ03QPWT8GDhs0AF36jo
N8lx6Dj8j1gZtRe97io0qkLKVskFg8y8ekYfsKWdEwakKgQBxAnAR+dmKdhlEVSw
oRmVyN2bmaTI1/sTs5B1qUd5q2vWwitfXWd3bFNRjUFnA3SFZf2fFc3LBdN5yBmv
Dt7RxK2z4G3gXWjwgzWF8xPtL5MWgoysPXIz7tXJxMXFCuLBcCgNNjRBLLBzJMCF
HyYq8U7UlKvs6hOza7z8sAnp90DycPOHf7qvv8KsLNFGSuWUNxz/H4sfEuL/NFG/
7SS8Qv6eQEHSQnvWKWyzM552RDkepWaVJKVlgcuKwBPKyGHSOEza54tXe3vlpANM
MAaqTDEqbkRPc9NPy8gMydU3d3h6KpLUM9W4g2mqvMTqxvOb6WA81477oQIvpr6U
8/6h5IE6wz96Hq37fj6GmlP8zTnL5EH0xX52rmAqbgKGknRBzI2042/kiGHlZUXb
1R7KMXvvICp1rRfxdWzXgjp/ciuDglUCvFqTmXMpvQZ79sDR+KSnWcQRvD/uZ2sP
7V7GHFGIEGiwRtWU+XSL8iTars+w6EOAjv9VO6YDg1wQRyTxq4VafuA7wrW8obU4
CwoyuqNDEyuZjOILwwGl817abbl+BBOqYFhULcbD1fX2UTRy1G7aGzn664Yt1cBj
uDd46HT8Dp/lJI7jLO6ptHGj9tY2/Q2PVaVh7NR/uWkbuxq82nH2ruu0qh0BZgMz
I/TiUiyzL/z8SvaX6X66GNAFIY7lCAu5MplTE2TF2rD4o336XhzAGoxJBwksIRw7
/Nmg3UKcmWAw4i0uEv8RplGJ2nXyoxuXO2frD0gxOj/MMt5E/7PAf7ri6lWpIe7u
sI32yIGtBn1Lt6m4Kpxs0d6iv1R9LfoYS0HZlRPh0kHyD9cSM++3rTAm7kFUp2MG
YpLxviJew1fLl8uWmpvLJnawlWGZ6lkRCZSKFYo/59TfQyx9Zg7OnZOOaJROZ86H
4wRXSUNEZUPJZbIjdt1azI1v0a69/T0JPCLiJ7AJvV70aWmthJfNOJy1ixiNHNdZ
HuXIjggYS/jcSW3zVk5pHzxYoXCL+5s5e5P/LSvhhwosUwQe5dnnrMEXetAOQN2m
P3zHeInFg/FbU3Wx0nCVfNWr9m49zck2iquaIudyrX+YwNcttCGolixNKt+UjSqO
Fi0mczHvXt4/HzkAvx0+TX0RjsI84FKgiLWltN+cpjvDrMXculo6YJjakHOM6IRj
kGcn2a5+fw3confKNMy8+KIZ3qrAUBRN1rRDTyPmlb+gdySKeyQq+qFCh7mUKH6C
LWK5vLdcdgIRw1m1Af9PhNGUb0LlyXDOTKgQMCrq5MZJvAs3fTJAARYJadsLfQU1
ttSIRS8MLqFHVr8mkYMzukqKbM4m9L8CVLiRq2FXi9TGq7+827m+YRp7qXt96NgD
O3+daRbwnTRxniNXJAqKw/x+33/eHLpiy2C7ZUHri/4yPCylGEjzAfzefvoOarvK
AVxGqiFlkyh368SsRfTSBkNQ6zq6K0flIdYahpzbJFe3sDF9M52VRmh/e5Ek8zka
kjdslcXO7btB9t0Aeud7XzVOSEJ9Rrj9QOMDzqaPQso1XkEoANQ6DNdbRLP8m472
/D5VzJzp9W1NekBdq9nzS4xPrjmq1nrVaDOCnzTNvN18RPgCwkmOr5xSXEB1iNN4
7n2QLei6M/HYic8AShA1LcoxPl8N8DmaD+NVU/MpoQm5hd1c2d6EiLUckc+txA73
O8RNO2t0o1DrWQG999PkjI6KQI0+HXDj6hhwtGIRD7/piaJOEjWfJ4KskdCxxWdy
rbmXiAu9cMC+IpEnz25VEHGD7XfmnbSh6aNe+yJ9bovyqACGAMm/wwLL91AglUnA
fDyfCJs1CvCV4+p1wJR3X10ZIbC02F/MEzZH6vbSOcsYyPhz+/k6jAVSzsnLp1vT
kEie6bQam5DnVHTjIZjaXIqoKFw4Mf4Xvb9DpXd3PeTrxZuPkNJJHFOgGmm0rVVZ
AK3fF7yIVn3mP7nglwxhTCMRmdxvbuaOce5ULWAIMq/QyAlUpJcww//M253y60v+
q2eRJv7dt5B0yd4hOqSypyShjMhJhHb616ZGlS5ylKKfnxexoRSfrdxA3R3xQr1E
FCGOhR2OgfhGG6CNsHtSr8y7d3SFJJ4HTfX1GiF9+6M9ZohzN7Z/rjFessFawxn9
L/s3mo30QybVUshXbUrtuBNWgNWaLzh+Lcr9xaWBeMbwpPnQkZYUXgxwt5xUy1H6
Or7t9FAO9DcKLP4V6pJZKBr/qfhy4bXwESgwWOxwtrrz6c3HJfMEHkf3FPkiYhEH
jiWHO6gUf3VxvDD5RuAxanUTAIQc5T3VyFoeG7rG58iy7blN6AOvwwyIe9r1+xHy
5KAyK3drpQQe9TqI8IfdurbSkjVoDd8wGjSGAVMxHHvVLoLt5m+HmBcM7cxFnW6Z
aCvaYoFlwqK5cAYp7dt4xsFY3l5nQ9R28blPQhm3M/H9u8UdmAuvXinEeIqwxOxg
kPpwBHqp+TIIdNfxYQcMpNhFAno7nj/kGY+B2CY3uuRHma7mLY5Xfs4yQ/yea8sw
iwvqZXwS+GHAoFNh2CchomsYy6jZtKHIybKc1///5nXxSeG8d79FqEc2ZG9uVCya
DumhKx/CIhAQDRI4d/Fkyg85zEMgs73MKgp/KzVWp/R4tUqJ7qzRRP3J33IWNJql
ObrP1jLR0jAMqwSJ1n7rUpHhfiBg8Bn3NiOYbaIIaC3A8ZBPaWiPx59GPaU3LHvL
n9JtQL+cSfWOH6lca1iof8B0++owcyVbPClWbJbZXZTqyZjYG4K5I1VQKPsV40CO
2MiKLQY8PfuRsiIjXFynhFzotpEnNPVe40iYxCItaP3QcVvaea/Du5AMfbvnOW7w
xYEM2LV6hUzi/FplZzg400nxg2b0F1mUjmhGbjga9lDXGjdCFTrB+hLDQm91Hd6Q
WHKUATCnbleDglKRApGydiByNlemkqbaKrG/hub6fO3ikjY2lCQZa+fqv66xs9w/
ot25jhClKN7XpahmPTcQAgtyjCCWhgcdU4SoJ6vWTGfvYbbNEy0DF8eRYDjG/Vb4
OtKmyfPFiLdxlphSDYZqk9zXwZtuDce42ZrlKqW2iTpNHJZOJk/G5JgC/+YExqWo
WxqADsqzVnOQ32ZvfzmaQ4NchoMyffI21fe8FElp5Q27zvlICA6Ut1QDQs/AkJJA
bpyhvdFz/jJ4TljjWO5JKQHFl060BWXI06ShVo6faKv+jQr7hERnbPgT3wGSoD2P
lY5a/sXHu+JcamFXQkEWeE8zpnRi5OvByNKHgOXwvkAwCniWKf7a+SU7CFWLJFNv
S2XsH+1jBFaxp6QbeGlWXTTZvy115MX/HovDWJ983w6tsS/0bD2rrGLCz6nhmTgz
pEYzFRVe6ZbqM1yqKHacoAGd6/qxH1AhmXlcx42Is2/gEi0I3WHhksaQr3gONaxX
WrboyCfbmhAdOnyuaTa4gpD8KB2O85/8qRmTdzUIqbRyYAAORBxW8tXdDd02oIdT
TR8ggck5l/Lgxq9iuHtkC7N+tF9oKtP96YtgMCnRzsfX/KVhIzcBmplTjxAWZNnV
AhFrwcrar6n9FHCL5n6HTh+Q3K2iGmAOhzhqowu5dfpQKv3/RASjPotAJRcz/HED
MoJk7mdJ/hOb2n9mITu1EO7HOL51xf9VDZkYAGvYCjQjpZIpfGTWdm6j0mQJL/47
roqP1KXq0fVIBA+R3VGUx7aBWK0YbHft6SJ0qdHRtcP4QrBU2Je7xDWrAsFNbSD9
RH1qobIhtav/s5nhzHEs/EyOhmD4X5CIfL14GCbkQkDCTdOUIbCzRJiswBPzL24G
1fwFOFC+P9KsgERteBnp/fgXze1iqL7b5CuxNtFNwTqGKEPeSAcsCuR2oXqHkj2D
bqIh6HEoD4KJHNvV5tgRE3v00mhOxpuzuGDAxieyFYHGq3V5M0zmSHpc3JVKxzTf
nrJrma5rtOgqtrywvty/f4VLj77uV8hNEGpzk38HH5otUqsNVKFvuZQTXffRB78N
jKZnhzd5lmTe+xdHUE2QCzzScSU8NnMj9ZxyO58q9r0NKfwMoyXL3sUGw45NSREw
lsMK1RP77nWYGuEu2ShtcP9lwdA3whI6VgE6TmamOh6e7BIWLkT8CI4lueTs56Ae
xxdhnW9Ej+6XLz8smRfCTyWS5Cccm5PIq+i18fQWtietOR3mzERIowYdyVYsz/kk
q4IKukZOjH9XrmkQnP/6PSbbyBofGprXpaiJ0yOLH7YOQWovR9emS61tLJyhERxM
PVLGhc4xEO1P66MqCZUgWtHE+JaFSyJTXT7CRWGPLdaabsfoqS3jW1qbksLfg+vD
+GmhmV7CkaAKEsXaVDpjr3XEMD2YS1OY0bbzmSCt/BFht+OkFJ7bke8bcB98N8ou
8mx6Di+tjnoTvYrn0MPcqXxZv1/Hlz7+Ckc0W+efsijieCJ4MPlHqTPBY++0Mh0s
qWPMW0TEGPjy3Q52VPph5JiMb4JwnIPPz2hbnZNdntnv/vFUylBtSpWUljnUMJO0
LvrQeE2vp/gIDaNmLF/RHkd6qeSQP6ZlBvZtafCMWNsX4VDUHyD7VfKi4lR3HmT9
TwXfIES52BTj1k1OfCnzaQoiM3o9xkJydNL6bNb2gwgykJu4J/jh04cmOVSekb4Q
0+dTW1mEGOwbLSmMCUi1YX5A5ZlguInHiaooehwqU77SRc//rpeLqV4Fly4BPMxV
cemewvPIWZ+XtxdxO/6/kFZAQQ7sUDo8ebtkIFCqQZu4yBumbh3Hhs/mGznGM5k4
fkdgrLAgjNZ9fCyH74wWGgZIHDZM8OO5x/Nw+FyFFYJpApx38nqfEuxAMJq7fG0m
tzkq4LfwRvBcPxPORKayzPDpDCFRj6IZZGn68QgysLoXXiTlZ0DgCBcZWPdc/xkK
WX5pMjHqp59A/A/F7G1HRw/fc4le++zpPEbWKubio64vwVbK0xbDjBKgtUPH+nz+
qt1XRP97wyJwoZ5A39pkdPthe9Ad9yJTIkeT0U05vDl9q+4oYyqB9PjT6kvOcEx3
tHuUpicI2Kh/K2OiSvJ7wgisUFuxhfnGx5c1zJZCM7rBVIITkLTqmCSKmpKPTQeW
O48XcmXYJLFzS8oTIQCWiOVJzq7sktq+benNxJwHs0dZnYLKNK9rFy0cYSyUmdVF
8Ho8GZGy6VW/f4TgDguJgxvqysNbbizzsarBea3l5M6M2U5fGE9UxMER8GHQCclT
3l4njMJj8yZg4XSJaM4liq4gFPPR/j0/nAVpNYqjwbdP/uxdOuNcKGBEg3RvWyEL
Hp+bjiK/9fvu2ZBvlQPPKjycZZbaJ6YgelHhE3N9fq9nW5uQiCmoL0e7hq/aPxgX
CogbOyUsijPlE8BNksK5okzmtxropK+0efAC3KUldlrBd+bU3sStixoTz6uTuIE/
lMIXMy01eD/gge45q4Mu7BHaMOQEMYHjXKOJj2ff+S4HjsZK7O57Em2Oq8JMJeL2
tiLYSnXl9ShAoXIfptNu16bs9NfIM4QNZDrql9bUGcvHjgoGXiaV4MAKZdJEXAa1
pzwNCjJvxtFProMGa6iF+DZSQi4ItUvrrbJTyHR2noHV4viQHrQk6o04DNnxPHUo
1fh9JO6aVqmzel6D1cEKYm6lN00857dZmoJ11QNnRy3XfZMuupFAYnlttr9y74P3
Olx5ls3gzH+E3iJy1NuV3OOJ5atv/eDXf0J2zOgxAnLnN41VEXsfmfP2uNqjm2nM
QCnBKemFWlxXwIYHbaVJzR2sZs/eAblt/O0zjv1Lw0PXTg2UuS0VO1mnesfzDvOe
m5ppTzU9zbizCNtoQdBbSXUFhmF67qIz2FGx6L4qPjmlkbQDO7rBJI9vmbby5cdM
7M9XUYqp0/CPrV5M9w1PHMKBwC2MrUOMm51MdWwF7h6pfFU+oNLBLeUyv4dFNhfU
bqIGAqnkmCDADl/b/3r/Yg0lJGS78xohI9HUDxjCnXbaVDlxRz4BoVr1Uz3PdCwz
q9e2rAcv98nC0SzatNCNfyKosFP+VQS+43k581Gp2SnhydtY+oRbnuynz2TIq1dp
Ifr9baLMOEacEG20S2iTSxxCmdGBuX2AYyimrajsZL7ODjCwhwplywf3HvI4zGsZ
xLtbQI+R2vkd7x4adg8EtYWHGH4Oa80SyPJOVH7gZTBMYuxOLqoZVyltY0FRjPQo
lUKKarii2eyyHMKM4SrVBVUYrkCidRvgfJ2b+GI7YAKFOZTP/B9NGZkXUa3Vchcv
kATcqDodNWsN/tfgDAkbbImMJv9cjMxn4ZxHN5WUHnaJsZQxUyekpJVtp5FavvHI
3q0VFF6k2xAIqR0myzRspC+Kq3TiRbLvU50ivAZuo8QuEuxouqmYgdNyXtlqVmu/
BNy8cwiXHM41J8tUxUReAOrkcs8ymSldPdQsFTg86gFA0kNgbe4bZ515KWBEwJv8
gEiHgWngsuTim9lyiT1wKfbTFroWgvUGLEo0ypSYKDL+E055v386YDEHcbM8KnI/
MogqDzNxHqruIsFnuUQkVmY7ILIex46Go3lE+iX2CvpZPeeyW9xGNaTbWdzgc4nV
ZlQI9nsW/vP1qhMs6MuZy2JvjccLmV33fQecTwobMx/0LIXttnot+vLaRV97Z9Kl
Vz0lfsX3GOiJV5Lm1R8KpzpGiWPImMAocYw37JUUoOL1VbtYBRUL8mDGuNP6XTri
iHyT7rc8GvXxlF5pDP3HWyLn08CIqbYQJ6klH+LRLuy4wvy/fyrkesv6pHDMPqoE
2nwZUlPtti2our+TUt1qAmHMlD3QmKS5Jc+f92zyQpidb3jh2pV9qSX04udxj85P
p6Wxqbn95fp5rclbExumwlafR4nVZhZGmHMKzxCzuihy+4oINlH8UQ643QcLNLuI
RDfOXZnK95Oaye1i1ZbgZDbnBMjiK8J5Zxjns9W/jV3ihptDaTmqsky9AcdLHTWG
n++Yj931mmhofLdGJPKg6hrloKF5HYPytDEoBIANLrj9l4E9nh8ARewZw7wI+Mrl
kH5eMXEPgfohtoWK1BJt7N7rxFHsvXRYx3JA5dl+l6ee5qWAD0isQ6yf0DKVq7V/
LGwF98SAXQ1pa1gMMPCD+cHLhA7GydU2glC9jm1WzUa6YfDP9xQGOTBpF4w8L786
qDOGgdxAwNM5wZ07MLAOk8hZEXFJYF5UtoKO8VlPXT6oEYVAHK+smTQ2Nrh+LeBy
Ny5LvM0SrycpUdJhtQIob8jvX5VAqlOyx54P0f52rvBclMTsalBqkaYIJjdfXfQv
rZnqdJ+7DHtv9WUPrjPEqP85LwL1RcsXvt04FRegIw/tVaYYFa4+I/Iav7s7ORTJ
GdZNM2CIORdFPPsyHUvHh94NFQPdatL5CjK6QJBJWOfv57VMmtyV96R81JZH+pCB
+GPm90Tzc6rbieixPiqOXG+/+F+A2LGpT6IoON2F3liTGqiGfCT+ppTKohURfbVF
JCYZlr1LY2675YXbXeH5aRHGZ7sQ+AgvueChpOehcqR+NCMmBUrfw3IpQ1NJjBxj
eFVe3jKHkQzOqv0VZGJk1lZdwC9vKwLlrB/WuVa1h7LcIQIFFT0zLw1wJDGHscVr
oOfcw8gHSRc/Kp3fts64rtXio9ZtDTuiDyzmeOnEho2RQQ0XQmYHNnyddyqyErLM
JENDL4LR9fnbHcz+JqSKvuu37elE/jUH4yjO1tccrH+ivxZW8S9lWlU054EiapwL
MsMown9sfVYhw1uZtXVFuJ3C+gC9JXK/Dpvk3oLtHXjfXD9ATxIt/YLdInK+Fzfj
CcA6NjVU4fQ//9XY23UYeHfw/8plnFNSBy/AIOntB1bRJsrReeovvJBNBGSXWQlC
dZgHYTbfAnS48+UgdyiPXNVmBFC5rfoOYI2KUVS7V9wHBgRbDcrqs/j0qEEZdwTi
1r5RzUKcoevqasM9SSPi4ho60pfTUaoU4ah8HEt4mFRlvxlttoKY34jJcXcTPn5G
pVYvIgr+d2j2jw8qTGqlHcNdRgaG8mfAtLt+6UmTs1jbBFR6nrdLwwqwFkKeRyGN
ebQgyQqXPRV4kln+7ZwiHxuVerLNCZwc5XK3KX9/NseoRFCZ5aYJYhITNj2nKe0f
AOOblQDtPHt7WizLZPDZkyo73Sp66yfzYMupqep1y0HGnbug6ydVQk+bBp35S0H4
6VwS3qw9JMHHDxE23GxemdrDL+9Nvht8PPGcoJs1xFTfdFvR4lSYDZzdyICH6c/v
bVY5PfBske4LBob/3FKrmo3vP+wTk60weeMHQ5K2DgvYWlH5pyw+TJ74Af4O3YJ2
meNCn2nIGLE+KBnEjY9EJJdiE4F+mjh4lLY5F/1XR6O2pVkcX+/gfO9XK8E1VGTO
x/pcNnupBN+9tEgfz4Qh+fv5rUoVO0BeTHr75wdzz5pXfxSVjIll7gd8zePid0sE
uusPmxKgEsstZeaAWi8Hc12WzDqsg8k9FJBZoeQu/1GVQieD2rdm7AsA7EhEI/Po
rWIbtLB2V3wNZs+54FgMPWyc/JAxsioJ1VjT4ATHoM54LGzEKiDy3FuydNVM28Sc
fXJSfPnMh0nJW5spkW4sUqnrgUya7fE8O3wdQXg4SDRgdxzOIFbjFp7aU1UurANF
hM7YEyDEoe6DOhW4MAmXsJJXhfAm7jfrMmtlPSFPb9NSJM+nXAUyCmFA34TIVqby
3RkU3YaIr90j7M3z+VvpnRuvuvIw3+jqikzwpoFo6CbkFZeiw9tNW4lK/wmloFCe
F/yjnvlJbEm/YzWU27HxFP8FcLHdrej4GKVbcjCNapFHH+6KqXQpmTokkQ4+qOp/
iCQ7VsC+3VpZLwqOrUYc4b8jgTEen0pfSCK4oKJiABUXH56MM7r8xb7RifBww/A0
54qtRzPKD0SHFzyB1rSg3Pu9GilHoZkiJyDfosVs/tmOZIXkJgzkDtbrtR7cyH/S
ph+wNrZXM4z8NhUrhJCPGElxGn8UrAbuYH6r7CMlk+AFv8FVYYszrFp2vi6gnbc/
3BuNdqwYO43sVBApFc6v1LqzFmzXoF0PcGHK5o/IWtSr6YHA2LehKq+wPp3RMuXd
tQ9lTW/SnGUpXrG6l8wXPZh2M8uCmneOvB9+/K8dEojQloYtM2lnSAy/GbgF1CmU
UF2k+FOUY84CgA6+7AhWiwRyZI5g6KqGC+GdQ0UvDJQDnw+0XUNMYKRyj08u3gEq
C/CRuBWDxkfDEKllVy0sKlyPlOEMRtdaKTxfhM0kBnhzWw4uFpCpzUj6vtbBTJPb
iyKfkGcQ+dHo0smsFlRJlF0Sp0MXoc9+EydNFxUYgyAJiiVTuE8lta2pixFkNmfl
gfMtomH0yMWOdsQelZ76mky3aKfvmWcOc+nGgVkm76ALnGPObeSvxt1rOm2pfdIk
TnC0lZS8ger/yKaXNI4P/gwFKn4cIkvMYK/SJGHKlJfgQE6oeqFP7HVyQtKw1iDl
lbPZm3k3YlTcmUMZu//XSlrZ+bt9vw9XRfUhY+SM03kgVLd0rchExPBuI9fCyCqp
Rv9CHUkeWlQbS38g4M60zYJtWTgVANRBrYLCeq+5NwvnrjPDLC3j4ojzc/bvqDDB
dUTOb1IP1UzZCcbh+u3m8R6GaSV8EpKaOw6XryVH7ZMv6vMSstGjYzXvUBVbnnxO
tTB4gNrHGgHB/4vmodJv6RbPr+IYRVN7CnTP1bn3kxsIIdLRJON7fPSDc0M/1P3f
aUSttLHhF5KnhaxyQVNgFIO59w9uUsb2p+BP4+I57cknG7bDkdJRV7KPwW95k2xz
/VPRmASF1MVaTBer88BCguqL1RzcKCWKNDwWEqeCaMiywxC0+I+oTbFetc77p6EP
3Lmk6ouRI8d/GvAY7u32a2vhMS/9knAQhtLmB6DWNNcMmTXqoJNrPBizlJaF5MIQ
ZmNPMVQ5LSrqxbB440YZfeH+X7SxnE0FP2R9MjYTBXDaKzkW7m96o9Nw7hwn5fjX
Dc9SJRZ6+gg046NVuadMpswkbCbchs/o6biZqfkRIJCB/xgeMlAqFY2oPJmuWU/9
8rEFnMvr4rL+0zYq3TdGwIJmreFmPodXRaE/vVm593Nc3/7JWQMSM+gi9kgDBaCt
KnSb+mmMjeFCfiQ/Nlt4ELUpTjH6ietWU7Iv+NCVWvDQg9p4MW9AXmeqrZVr99qG
oiQgyqj2qjk40hkAmYkIinuTNs5wwrJRvsZRaCPrzQrIzs1jkkCQiQnso1UlaSNP
jiamTuB3EAst8Ms4OV75zAH1jscVuUyMuQYmHxUgWOzI8idADAaEmAmwV+eTcade
1NNaxEkg3hhEIigRIeaAigdu0h55a6baUwiQAhwUYnMZij6y2nP8N2A45X2oxerb
+8aKOHjbeQ2Zi/Q1bPIaf8v/Wr0FO29Tyq8fWJRSiCuj6trHfwawn2QDLZ8Ho41E
YPNieTV5Bv2uycMfki2xCuuQTm5x61xoC+SaPny0BagKIMLQ6Sfc/Ncv3Nh2oxqi
v7GlbXqUPzvMpl2w3aoD6D+Rebfw3RKM8dJvoZSLy0HvDjh8xTHNEHEa1u/GextU
g1f3lwYJksR6OAumI4KBiICLGv2GmPj2B2ONVhd9Bq4wj+OK4la854X43OMC9y0f
6Kfv3+yAz1/Ff3MUmy7SBzXKEg2d6vA3Lnhf+yHKV04Ecez2lj6lNMR5AG5NKZRO
lE1t1TidaGlxwMiFeDidkUlm+Z/JTteEa/TF/3vKG2FTZRtmD5PDkrxgb9PeMEkE
860uDPyCaUCHiX+KoketWTP1lD14qjW1wSJghU7/2Lw/5f/MzLoLXiNw3Pl0IWKw
KG4f0gNcesCyM0eSmZ7GW/DHnGnUebZFIQJIaOEoOgjGdeReO6nIPpZ/ncYhsUqy
ifg6//5oMlf91p6zfxEi6chM3Cg0gcFWBfCCV69bDCAuMrte3nb3rSdAZta2QcdZ
infW0YMd/PN0zDXg/JZI8spN6veX2ff2CTPQcghJdqSoPhkxCd9UaNS3vqidl3Dn
F6IE+bq6vLjbGLKAVsJL645Dx2hXLZypmtQvqpuI2iYLsCj9Spv1Tsxc/WY1uxG2
LtnquDyGL32ZYuFl5VINqLYB1e2EKEDZvuEiyDrDxCva8ouBeYtGRRTfaJ2hEMIe
On/VnaxOEaHKb56O8ATd6xteszDwobSvcqJlZ3/jSBzMaBINOjhpWH9gMba8bf2L
LqDfy3cZroIZeXBrC7lyhXlRvNYKSM9bO4Bgu8UzJc+X6rJbDBmFzTsaKsOJr+Uu
kglx2VSOWmkWLJ7qwLeGiuDxM7P1dGpH4/IbdfjnW/hf5j45yTU4gKQxJeomBZtb
PqGOvQR6bkN0tc+Fhn/lDDeICzw14SfPsuqwZq05K/h8nhUEthcFCedqDMpOnV1o
TeK1vnW29oYGEuNTrBzZKBP6CUdT4E8EZE1er9nOrmn7ig5FM/N1nNfcjz/Iadqm
hyoZdAoQVPvNSGl4kzRRikAeoD/B8/R9CbLhrfhOhT71qpUr0yKUDZIOuBB4Jh10
5rVFiQTeDgmulKYFd1JEf0HwNJrCLT0y2TdHo5a0IIkmceODtyvekmP3GFKM5TGl
qRrRECCoiBCxRRLiZ4G1JrHSGPE5W7t7DYGlTqt3W2Fp7ZgWjrbnZcivGU1PH5+4
c0/FIaIg3C7A9dd2nR7JCuARp6EJsUCkI5glrDB3zxetCrizYsV0Tz8ix1euqspw
BYpoLbSwAzzWGiauDcuQ+cxVmukHcEdYY+BeFkfge+gUXXB+jsMcrjY85AU8fr/0
24I+ZUxNb/Ycma07+wI5TNLCaaNWD8iHwwZCbekscvXSkt+akeKdmXlrR1TlUlXC
QccRbehFSKiI+rqU4alb9zdX2FjIec8H5unozwXRoWQUDwsfaod9SBKJIBJixyTw
QrvygPhA9MvCAaNU/HGozG4gmkg8cVGtKxnb/jTd1vmxA+Wsg0LZxc2calLCccpi
mWiRJJQHC5WLew+OQ5M9dbGc4vSxDOdBQSA4AgDAV3aRwlYMfOLZ0mwYyX5SLRUB
MuwJo9hklxarP64F+f825fyFVfVJOrbk4M1ect8Uw/U166v3nlvHaJta7EV0FIF6
eABJgxrgbYSsySgIWl3jfBzUWt7Z1k33WLUz6TEds8J7AEA7EcNPffglx5tf7Y6o
rQ5JJg9UDva1K9r9UmoEIrvCaD35Zi02hRiAck2i/zyq7y3fQ1mZl7xZOkzifsiy
W6FgmEXIfHdave/J9EmKGJ0Joz0SYU69XC0BDS7uyDQ73CJArMKj22XjOGG2ri25
GhxtChdm+rPHLTmXVPpDTAxSN0dsaObcSviv3tLJC5IW0tpVfWNbpCUz9335Dkj5
hGCXVYQ0JwOD6h0pIDczDmvrV8yAsCoYS3uh2J9+/oLuMrLpUssXYEK6/VGU7IF+
TFTyjR+3CU0bszduyEKtVZsDLcG4/MHLTpw04SsvMcLNDTanf/wxp1gKnV+1Vy2i
H+bcQL8rT4rD1+n46LEKKnR7PgQYlzqlF6pclpI/UYm/fHqxRkFmSzY3SisqRP5b
Ix7/04POMbfTE7N+gIPQm9sRbJq3XlPmk5dZnBSApZz3AGQ6207izgx6JIt6Pjxe
Fm0hYV6fX5+FFiEAqHFxrGKeR3VzHPlLNSDnqcavKkox0H6+JNrQnjJjvlqziq6f
R7iNYokCdnjUihNk8JnCHZ/n0Mv864ETvpXpS71n+wBC73044OotTwKYhqzVPpi8
0dXDSdYvRqAaEPh0kSWX5SuOegOBzvdhpPmcmq9D80gibqpgu1wR2BtygXuYkEPk
bSsjCU2J7b4lCvsBUFeQ45P5wzSiFDfLQJeLQCJe8qDWNVIx8okBBgEYU3yua02f
h79+UeMFAZc4vQFy70zxdy9BY0XEhEFYgppQ0jEvT2+CMw/G/qOLN0guiDmMtuXF
+7DS4+PisE2UuB4RMSRaw+sUNSAGF6tlekbzhpfzm/Hc3PiTDw1kGujgmGAWmw8d
HZAs7DJkBjJ+sqcQzbOqhbqgvFMeIp6WU2OpF39sCB6+pS+uVwFHrc63cmCGF0gm
4DHGWaifOtEov/18jqBZPiMmPVv/MWid3suHiDnv1vul8cJl8fuWSdzA85Uu7ze/
WlghpQKsttNlSKjTuxQm60dw1PqwQ0ulJxr3Wa254DSASFd4UIDShPm+a+o9ftIv
wC9haVmzWgJzQabu1+u62DSDkf5r5DCxM59XIH1Y46E6/zu2KTUxBs0DxXPrBquO
8MmOVDpDM6QBxuBGe8PFTCT5gNBzc4p2dtyy1+6rMjhoXBa1gYx830XHID+vebkt
Dz3k4XXW3cedbVsCPvlehSfeNR8vIZ9BBFHQoxPEXlFuzWkzsJcJcHhNDs5d/TQF
+pzMb9+TSQrufZKE1G24A4ILdJslcgU0FTCRKq4g/E1mWNZnRXkcHkj/8krlzFN0
lMmuSoNd/I3J305v38iFdibBsnxCB6VI9/RysOJwSvCpYlAmFXg2KwWrP4aGykqw
upCFVZNTcBSIkTcm5ywtAs6VXCQhE9qwdCBako26HumHvkaSNsMXaSIqnyGH+3wy
MYD2Meqbg+Hdt4Ox+Z5UTakj1iQpk8F0sM1bPawF8GM+EXv3lqsZQh2V5YT8fGv4
A7kIp04J4kuCNLYEY8Mq7Apnr65mxvdxJXXk4wtfeSIy1EFN4rrRnYFOXA7KTdb+
jpF8XFZKtb1svedZeAKCWtZ/OJ4zH/6V1mqNxhPvdCU6kyvy4ansHIHVH/IpeYNs
terfxKGNFt1/uLiAqydjY+uCuWb6JR4gQ3Yi/odTmBlZat5cf1Fix/cj0O5iW2Yg
NsRYtsPSk1HJmL5e6Ld3BZn9MdxaR0T5Bo5NuTR7sJnN5w9e/GjKM1tWYtvv33tL
ft0X2CK5BjI2XqJs8I1xEtlU14GiV/OhrK9EE9Fhn3HfUe5BSYWyxKwWdyGBfAuI
Jr8FLlinkBhdfohbrmvOik3NHqhHivIYNunQwArTMkIPKMYkxKogC3kodHsZ+rPZ
+pz4KEIdTXfoek3QjL4fIsls9vJTiFx5tWjtIiAz00VYaMT62iCTcSPmWxPRYKfl
iklL9zCRkvP31hoJ0D667rJ1713XRWbCt10ETyw0kW1w1njHuSnQKmfMNEGurRUw
uK/W9bpqqKBzNoU45TB+9FkEnt3/nu30wvd7OuuTpznwHoDdoBG/5Qksuko16rIe
459jBp7r4ngLQtm+YOauCoUcQU0PN2yXmBRnYIV8b0CFtReYQWY1+eoum25Lw3/0
Z+qme88ev8AvEA5Yn+YvKcXT+MjYdZxNU9aicxV8Vv4HGc1x8mShmbOmegE/LyML
ElQhMyXarrxrqe/2Tazd0wQ2Gy7GrTFquhejqN550Z8qPJp+RUNNn6oZVu0+d9ww
k3ZqmttpLhmLgA51LuQB9ULZ2W+T9M+ak/DZZg9AsglXlhAUrNHdTPO6A/uqcbwQ
F7xVw9w9LAsEl4pGwg8R16F6zEUvU0lW41IMGUoFD+9Biu8Qw7IU0a1Ho1PuSDq6
3KbL2yUgeir/DdLA5RzP9b673AQvAADQEGeyKlhPBaS73lclXPFWEDRfSvZfFn7Y
v3n+EUSEski6E1De6KIA7Cwyt8Ah13wfBH2Pw7mxOTPn5gISvj2tOaF6xSa4TAHL
vPui251FWNN59iOiZ1WT+1c6+ywdK6No3ElZlEq/rpWYIbfUwzjOudqaa6cISBop
wYrdZA0EpE9gAoXb5fQsowAdr8KIjUNO+bwvJUTUHBHgXfyrDs1xzY6uo0Bp3iTi
olxq7ygj8uNUgTxqavnKarqamIGFltPGp9/BlfbKmr6/wnROmHlwS9cg4KvsqJ++
pe46HjUAQiov9uUzUJV24fG5gSgNwoU8aAAGBvWEbRKZDrWnSkKAY6AxtDGXg0wN
u9ci1Sica/G6dbIXEgsH1girRSJRW7kYQmmDOwHJ26HhZ8sOU66Y5F0BEUklfEPS
dYONKd1iPJybWVNTR93uZ1OBIR8NYcG06aEHqsXvmKOF8q58VFlPfQRgO/Z3f/yk
gzwdc4VDa52QACNLVZly9J+7glTxie2+9lt+iMOFK8fYE06XhY4hvqOruEGu3H+D
SflD/EiIRMeJ4UDjJxAlCA==
`protect end_protected