`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10368 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
YachDS4bpHRDzLXFQC4CtbN8lxqE6WQo935aAH5tNg9sXe8hlnGamiDuJeXoNnfR
NZABoaTI+C9BXZWRzAVE4gfP5fhVwHNRU3DLjPZk1noXtt/8gMukmQ+FIKG4XCYD
70qss9grSeQB28Rs20N1yamBpGt1W0eenOiRBAZCATRuYmyhgoqWr8R+jCh3c325
n0ir4XQeh+4WkCX/x6QOTVC4RHmTOBk3t1rqytRHwjuKplhsJIVXI6jIaY3wrw/C
XDekXWvQ3sj0usyeK8Tj6Xdi71YKNiktgRjLb7VJayUBcXBeTw6ooVGLPF6GZDlM
mpi6UO2oeHQvJrVNjrWz2/cc5mdhzd/kTreHoCXSkIhkSFqLj6pZo1aOxehxFDlh
RdwWKnEv/kW49nsPKGw3aHque+EAuAvXRIetYSdT4fBgbDAOKPTA2KJbZveOfhec
62sMtc+SriXMLgpOOkLKkoDFy2JxIzTON0oOidvfBP39oR+h9YfpFCbgeqhOvTU4
QvfHgbyFkBIz5FqNStz20FgPaib/+Nsqr5zog0rd+c/BiOhKJgriCN297sI2bEXK
Saha3zsQAvG63Uhm5Ve84l+xgDoWoHe3Giu2YU5jJ56b2ZTvx+fvlmBKQl4JmbqQ
dwHVLZhrC/L2Qo6tnrw+jSi5w2uIxTA1pHjSKVTado0SYmyRkRN30CQ2htZc4e46
1TVn9nul40H1DJawiJtMzEu+1jidc4hHHQoOHhYmXzWpNAIs/MkI2FlPEO7G/8O6
lCdX1BnOol8OSuiacOALHDBWaYHB3QVWrsc18k9zMo7WNHep/IuhSbwZ0n6wDvot
F+jmPlfb1KGBGDuSTgu9H0tcyLjFIOoMcIocAN2BHQJlTjl/xlO9fBzBQK03xQuX
D5h97RjIq0c7uho3oY80VV0EU+QQh5MI4ALb+GX3KTPIMTGgGRF3+gW1aJPipMiD
tmBYNfHew3/aijHVN2dG7f37kLV+tETc14bWwJvptBfZcUyqvfZElfb5xw4VTE/F
NQ9tgEUZt9jX333FCXREEBDJgusUI55JfPrqAL8JXM+1ux5WkVbU/nkkyWdZ5+jN
Zahcgma2J66DRVbejMgtIRT4o7ov3QrAbyF1AbP7//z8C7POl3Tsu6b+pgnyZfgI
5YqC722Pfzn5AdoyTqmO5TcFmqJQGvDulbonCNyFfTMC5qtrqOJCKpdJdXTO6Eef
sal6HbqSOS0OJ906eprhcFWz2ocPzKw+QLBDDjqAITu7gmaiWFybohe88JjijHPY
3pouUe/sI2yWFhbV6vdhuoa1hyo85EKqW9vFvlaLPRwsiRdIa80CsPbvSxG2e4Zw
h7X7IAKEFDQudqqGfHjauoM4VHaXWrsSv7Ybg+/SSnPF9Pm7nlERitgoces30NEB
4G4CN1tBeC/AHAL5Jk/4EwsnQxp8NM6NbdoTsJE2iJ8ChZhTOPfONDPXs8SEzhct
e0R1DpEQ/ksfpYe7dMkHbvMSTgZ4uTpyStvFIW88W78uy3SdN9s9kn5S+px/wenc
+TJwCmLJGjEbOXh9TJRjxabCPjII1ao4v5ALXS0ccqBEJN+ui1HKUUBeWbggSepX
B2m0GYqT5Ngm5oLjbSzljeZuBEi6vE/Jk7lJfsc3MR/jN3VxFOQO+a64JKZgVK+q
jgeqSoQ6BKcKVYvUzNkeJdosgz+X9f8e996LrQVcFVlyGICwANfaLRHyxq7Cv638
3YJEe18x9mjKtSW8LA/UpN1neMx08fJLDkUYWxg//kINoOzyERzhE50UO8az9qgO
0PlgaEfDOzS5VkhsmRtaz6EU0K1ZGHdLoCp9jPs8/0jqQFHPgbStGydQKx5K+SpU
uIYjGxzJ5hkH8xXN0FclC87jcEI+L6qBQ5a5lpa9pOAuFs3vu6RQxFcFa+u141GH
IUhnCJ45cPBXYdtgW/qA3+IH4bf5J48PCNy1saSWRBSMzFDsN9T4KFoHOquHQb/O
bOMWu0j3fJduk++BovBTn43hT76cyPf0HUzSR1k0xaau1rKEjfXFIVv7IJ+aUOqQ
Y6qCzzTXYMDWSyXlh4q+7cQjoURgVJlpv30OGRqsCBnXZG43SZjuPy7ycqfQQ5hT
oxCExqCy9P6zSXK7Qp164afLXCe5dB9fvE7tFrIuR3nSZm2cp6GWYY/OxABNTsi8
h7c8Kbk6oHiS4srO0lWQm4X+3cnxpOPSzKBdKcAPOieMdX9e7Ha06yPqcD6vZkRr
cAwKmC0yk5ArEkGYQVNmt+LlepTlwjGWbFMTAVF3dBCiRd/1X/aP718i1auAyz1y
Pl2XSw/9OTtSftFlKQR5Pfx8FzkFnd3LCCog3z5gNa++dr7xKFNmhhmbnI2sJh6v
MQhMV63VvXFysE17f6niyKw336L1db4IxVciHeRqd04bSiZL8OJNjM441AKzc8Zd
5iyBn70z+Ayh3EHwJltkEzB59omLeFabrwfGhq6jP50IHWoxZYBnQ9xx23kpMcvX
5LMH5uXtgYcGcWc9EprERFVg2uoCJxFQ//gpge/V5XIT/ijtb7IP/WgHe8sYgIHM
e3rZgmQZYnGzfxS5X1U+9G9546yZxzLp1iOXD+SzMtdlNhOPpDBFgzx/cLWzfzgu
H2OvALdVbpL4It/tOXDyMKQ27Tn7RWBWCE0bhff/MSnzlnqgFQT2m5wC2HpNqJC9
xlalC/3bWiBoSrJysS0VIw7UcddvA6aqrPByvx4ODp4lnxoLCfQBUQdJ8829enoQ
6JOJ4Ph9jpmkGRe0ul2r0hRtlwuK2nb+/mp7tmG77ZHJt5BA8MOaExjOkSOtT9hU
RvEVG+8qY/DJlUPeMLyEtgMbgKH+gUfRfWQ8hiLkv1BQYMyBjtKfbdouRdXWI1Br
odW+p9gWHjS+kjkyTIwb96NGv41WpxxJiglB++rb8b2f6Vrz3IKRTug0/EXnk+Tg
WHOzGOv4gkL4Y2ugKDhpXM6Vi0k1tUueToViF3QxHcj3ae3JcL5oNuKBS8vtpYBP
EG6mjUu1yrwqfjheVAUW2fPGVUTV8Omqoszgyx93Ae/W8fvdfRXTyXXlf09s62Ui
N5mZS2Dcvihqdyfv8pWcijk0ZSxaGtejbrbqQLaGRxtVBNDQlEVeGfXKgKolCc9I
rhzZ5sOVgovgbnEbC/GxR9FtmeFOMsUarNbKAqkv9GC7PGiPWLi9rTrdDO5OlNas
MynuV6KNxT5rYLh2GI/QGuGL8qn68EegohqQ/tGsOLZfOfSoolVN8OZI2UvTcwyH
bWX9E5J6X3vkieG+TptJOdm6iiEHTIAr/qUd4Gnma/9zGIWE0qfLoVi51Vla/bGT
COHiH9Ju7QgQJMrxDekbDgd/ijpIiwf87U61A5/ntB5x1wNj70UTsXrE1PADj3DK
8wGHbtIGa+rjLi4UcMVqe/xlPa3DjkvoN2aPe14xz7Fhjk8aNX4NgWUFSJpYJOKr
mULn++feu4JNUZk95J3y6Gntwbi72K6q3yvneWuuyg7mNmmvHLCCO13xKdhJvKoB
CVmwup1msdG+VzO1UCQlqy4H39Fw431liDjoYw94kgyJy7zctSgZMN7T/YDDPt5f
IQs6KUipRMDA5qeZ/wxQKSedUu9wteoHnDO/TGz4g9+NeyzcP0ImD0Lfm3OX6B2I
F+GZiju27Me2hPgluKQ5whQmwx9nI4aykRqgFCLJICN6hdj+eva+vPm0sQj/Prnp
hGhWnjymua5YAYKhtMYFrngKb6dl9fDHmYqPDHPdNqhFVaPjPikl2Web0PL9Ru22
ShTZtFWtZDyYdOdx01M9cdPzzdK3aQTyKIairs5YHk1ss5k+lwHUXJ1yWQJG9z6q
SBTm5L+iCuDMaB+LaI+FKxS98115+em5BkLpZ4ToZyEF/W0u2vPpTIGrnFvoG1//
5XU7V1Y3NIEHxT7hBMTrLhIDrIpqbLZNRahy+KmAqau50ZhFqpZjZkaUN5fTwMjW
dQ7/wy/SbsPRYk+Py4/rdt3TMHuUk6tsiqfYxI/0ZOiMYuZ/H0ZcFC2IGYiyEIU3
gI+4J4LR0BTQ3pFnar6uWbUBh1cpAeBoZqd0m6ewd2Cz+sKYnkVcMv/iNjTh4ipv
fdk6Vap+Ith1ZWjB/PXrvSDPSv5cyHcndMITQhb2k/NPALZJko4A/5sNpp+bq8WL
gPqtrUDka2+ldVdfyFfgeBqHIyoxz6wR45HcoFryVeCxu6r9bkpQ2nRrHPkN8L9I
0698OiIda1oRso+3S7S7cBp14MOcz4Poqxlh9+DXMEkTJE6rlgyxl5MN0xZx7NeT
ABJ0x7fALAR74TXn2wG3sCfzKAHgCw/SUXMsTg0NUj6Ie2ieVgcWQdYJNB+B/ST7
OA7udHjhbNhtwQQVfPmzFGPY3EB2FBe0o9V4Wi1k/SGWSr3MNjfW37ziRtKPFJKa
A3nSw0HBgE+f7ykaZCm+87zTpEDU0a0vdZfq1W7HDbbQ2Qb0nS27vnWq31jPl15X
Lma7ULTCwmzLXGOiWqP7oxa1e5YOslyEgF4ngYmLZU8H9cov8yNP4YeM0M+St5bF
i9qOhyZJyAScFJcaBgV8L08Nmp8lg0VxWV5Wd81alv+uj/HrMpkGCqcycfUPrF+Q
cMGYJxUP1T3nR+MeuwWYPFbvY4zqFF2/STsSiRwxwZX3kGonNGVF3JJxSvN6vLFy
ekndwAqJQ/PAccGQ4/0E7QMJ9dbc94AMMfdfTM/9/bjVGQ+D2luKztsB7FJF3Ff8
ZL0PWaDo0rC9GMIFDJGkAl1neCx/z73GlbJ6HnwTkVC0nIUx6HDMRnZ7vqW8TBcm
xMiyEte9YedpbpOB44vWxBOQ8fkYwI3wQq6UpRrcNLR7yYecCRzH0cr/g45lCp/2
fQbSdCsInBAjRwQAlrv0z9EGWHS7hQ0iR2RHtNpN0hDVHycy7QIhL3dwpEaaNGUl
mf6WXQiPJhljTkowK/G56hAVDBklaODa5D/v/hI6V27r/t220bYnt2UnKLWjklO2
yCiLdcETOYklq9lHUrVwNQBhGkrq8fnkJpiYRg1dIobn57lyqtsNPwTXiSSPvmbX
JM9XiXl4g91pZPdVv+Wuq1W0knN7MNT17tw64oik//MNMRoRWREEEJp9XDT83m/l
CJcelhS3aA8lJ929+XMf4izZcJeTgF+3GFePZgCH8d2ESnxsHXSMJr+8Px3N/rGs
nW25+KoJvRY0jhATOX23Esec3qtlTz/MhDTo0tp7bz6vtFU5CXx5PgmzLoN2PJVJ
kS+B9+0uv77GBIcUYrLdrm/k6pPxD/ApUl2wq/+6cf2y7MD+Q7CC+u+HCzUiG18g
nKgBbr+RMRU7JE8VQ/FUSD8smRvxqZ9/PEnNbpIBWgOrPzIeAsrEybusAURqTixg
V4rAC5Ah2+EXH14oteqVlWEoNO+g3AL1cK+8S4y8n+skhhh28bDLx81/EYpdteBj
besEAbAujvPmKeoKyx+R6/Nh5L+XnWm+W2voqLUE0s7G4R+dwhYpIvBcI7hbRdxs
7x0xrr5RCTIGNbNJfy6sMyRGigm/DrVutQiC1RJWWm9aPBx01RCurVuxNSKd8qFM
figXuZXfMmTXrr0WCu6f14PGZ6PqKJBaKUdEeEeoWSiEzWqBOnYGuR+27RWwB5Qv
/U+DijaLNe0/7S1v1l0n6GgN0aoKRSh96IPyUYK1zx0Y/p2xNLmHndxWPDsf+e8u
kSN5pjugDZnjKZqzp1bDHxQ/pYL6cJkuV/hlZhYivP1Qf+1lRNKMDJEDcDx5A4ws
6ZSJl2PLoLEyPg6lVnOmc/z+9btsdWRNfkpDNYbX3b+1p5SR69TuwJhWzj3KRu+2
hHVk84s1rodskxJrPrgCvXSfBt6lwKD3/Jbj8IZNGiT+NK/9OLhVovH9J2wk/Bko
A3j1bb6Mi3I+9bhzKyf8UHGUdCqN4jyFM4O2gxtmPfvt0UvWqyFsGnHWlR4p7hid
2VJYMb7XDq4Vejs9GO4N/I5Pj26HauNcY8JjG3fyJtNwyD7dX4TdVBobfYA4MbOq
8ldE2+M1TVZz6qcxPwl3VygQ0AWON0iCAO2xbwpWYF9ZAgvaXkm1xcLKQdquBJ4I
sKA5VAFRGy18j+mO+v7nlHQRBtma/8kPDiedieF4GiB7gZmlqY4Om/KfbjKh4nts
BBeAfSDN3d5oETU+G76vTj5GlVe4kNDz0nCaArIbujCEVNezH3dhIva518HXG/pE
Emf58PdP2tXvfy9ypHEUbGD04oFaHej/uxiNfjyKaMzR2JUxXGjKKsBmB4jIYrqn
0WyBUHLphoA9ZsSNYXKTk4CsTQl88FWT7DawaQkRU8SozS5rnP+UMJWGWrA+4lai
n5K0a6utpLESP1ujTNTmCG4NYTFwiVNmzYB/gc86RlAB17hOqonne9Bf8cbwaI61
8kLyPuRZUVd44KMaYVvaLvnU35RyhwASVqjkNtpyi7XYDgJ3kWKBVutbrhvDmtmJ
jnEEVpGy/fwJ36uIloAsNoOs+9UofrQvQTIlqOP0O0CJf9Mljsv8r1OL2GfESWjq
pU4EB0y9ekDLlMukedfnDuLU32UMCXNe1WlE6XotGFL6o/f77LjrlgRTqO8XjPqv
UolHNSlgJpC6lLDh152vwOkbZCWHh2Twf9jcGt/3OvNxXNAcMy+QKPJq2zDJvT0Q
2tI/iWdksfDqMreuw27/5vLRlDXaU7TOWXby4iXfSqD+IlQOvS1dMPN8pbAlCpxE
jjFtbfhk21c/TSYNdyMNnh+C1gn14HTTQhgaNAbbHQc+6GZkfNa90ygpOTIfL46+
2Cb+TPzoyS4yCnKjV95y9pg7Z9Pe42S7+beI9DJ5QiuTHvrnSS2s8IOk9Ibc8WCK
dYrc6BOix5atTxOUGg8s1Drwyazrrl7O6d+j91H1gsUf5RBN14h+efkzM7Lr3Yo2
At9FJWdujImlQDqedW4JGHI+Yk03yHvwyzO08YTyw2mUgHLxQnD1M+v+KvTbsWrC
J0v9lIfXJJ9Sd6Gr6FwJQfkFUC9tEs46c4H9wNSEeEWTvyKyVadtLADBMjQpGVij
EfoMWlwW+4nliK3kJy5xOUCXGk77tzuf7wU4YewdpfYasBUnS/FYjqkaU9/AxOVV
BhLGCHUp02NMG+68DyoarNdPH0nwxAMLLNVriAU0OFQV+9aW5UiZxgGk6QttHOUc
xupVa4+Uk8rHpW6Bn/ffJlbKT+Dc0uzysReJonSNzjPEqBOGsbIZvmfcpQmA811F
eqW89OGKhA7odyyfSHkTxMa9Akio6P+cyx2kUCOdnNm7Qp2L4fla5+YDbrg0ALX3
wuNxYzF8P08YOmGHD9Hfz22yNzNxO/9kWBfPO+vVSyp737AQK6oCn6cCVGfGna9/
JDvjrE6dFPqg5Sry7CI/eAJYN5Nw2aRLxvKQTF/eoKtIEbOWubqJlKSQIjzDa/ay
vo6aHPDuF3+unXNzwtTyQpNGbTsLXmgXXmkkynRmgpJH1K8/oEE8v2bWrAzUFXeV
OBLcNfvImqA59KbUp9NOPzth6AVTKuaTtxZ3PYGtZJ4mYGq4NkLF1oAb6GFNaX0E
inT11v4PmVVB6DR7BG9pKosTwO93jDlB2me56s6jn30c65gIh7IZFwgXu+3/9t9t
iEUEGk4J5RDOpxgnDmels7hr70FBAJz3m1RkJazhp9W3x8YR1jB3EbwKgMRWbUhc
I/hOOHPCOGMJAXmam2qTEI1iNJ3AKtMUUEYVfr3qDEH0x644K+bsS4JHKVd7qehF
Xp4FKh1nkCxXpcBh6aoSIn4aSVXPNEIVvqVx2QUGP5CBnFyA7DBF5NYbrpF5BeyZ
XfBeMVpxmwA0y7HQa9Uyz3LVv44TuDW64sEeZUSj+ZeghCOrTjvobzYCgkdh7O1V
A7s3xh/8W4lEKX0uwsbaSWa9DWMGyiC56XUPnLwlDZB8Ok5w/ePcyJSd3mWvy1qQ
AhW7xg8n7CQuVbiqSKy1EStHL1q8N2bz+WtmbJ+85Sb1+DHWRaMA/o+n7FyVolTw
v1FLQK6VtYeVyf9au7BlULg/jEPIKsjB7Ezo+nPyP6DJ6OiAXPZUINbXMUEgUsZQ
1aUhDmJJLLq0ER8HOWpsTo6HKUQdhH45Kn0zYbQFNrJJ/cXKqgdBPGV1R2IvRxFz
kTfffn+trZ+D3hRROTsSl6iaM41gOkaBsfh4g1g3TD+BXkxdzPAa07ebkd50IhLt
nSVGJZ2ne4Au4/K1SWGU8BQ1uSn93yHKfzFrALag6CrXD8wC/sDYONMzVQH+hSHI
JdAAj58JI1exLddq3LVwZtUwduZE9VB6jlbcW7SEZHS6JAw+Ga0MoEzGjjRdrFk5
d2oWwc1z2wJRYTRWdG4uEL4oPBoK4CKvkBKhac8FF1bd1R58rXgiLIcGfLOkpWnj
e+HSYrM4YXaqBGh43BzgcBgzY/uWuRuavHCSYj+SHQrGyoIr3fmPQPw7vtorRCxi
vGbN0lK87r/EN8KkAWMz/hLoeDuGSwhwXNgd8FvmfjjhzTOR6vidwPzWuBo9czDJ
NMCKk9zLTxxV1NJ+1hDDDeamlBhzcNOoTpwSp5X9RdZGGRII+hyofDNUx46vletf
DQTimFlOQ1RbldzXpmfjnTiCY6dzgPCW5yiqWaLTuh58ocw8/uKhQrGus3wQtAye
aMDWzbrREpCVFtWP9AIsw2in+7tP65WNeDS2c/upWaxMADh/HwgM0Mypjkourfo3
y+1KYploOrkCwu80mR5ETSRTmCwZV27ijn/mOYi1nnTmFHAxxZdrjapEG+4SSgQf
RsoMliw1yyU1DvaJp5mS2M78NdGWxaffr6vqK93pGZXOo5d0Gs44O3Bl9y/NTbOy
XWoFzookCEjSGo5/wBp0I8/Mjl50WzeTr6EW6W43JSFJ6VkIMELzfyHZZvxYlXnz
vdCnsXmv/mqI50jXo8F6pPjpGGuNoGb/oxrsTpfrXlrOrh8AmsPD08W0NR0J4CsU
t7B7cfO9PqJLrcXnvNuxeVrCjtiZ4oItpaWtpjZ54SvN+vaGlDPmyFF90Y7yb7lI
I5m1k8hgwNBnXTJtmHPUSQcL/cn6QMHerUDdoPjzgMt0L8aycHimHSboDT56Y6dC
SIwjzfgbRgLlTjTCjaiw/A2B8F/guU047XhFxSBH2pVNF+bXkxCoGrpvy9Bc2VQ/
aZvl4g9fZGkjjqfFa4cNMhm69T63Dj93JIBhieoiUTHG1HiHDfRlTsEE8iRgeyeW
00uG2PL74XCGGfJcE+xfOIFSEf3g1AC5bTQcWkkkSyi4qj/ekDF01ZiTQ1zug0Zq
sIAFUEX8ji7Xy123bOpAf5q7ITRhmPqcp62g73r8Ye+HfrHbKjULakPfSw62WASa
hsGbjGn+2zNUDFZ4jReTxWQp57AoyOi0EbqJYl7LchBgeDtv6NiapRHDNBx33nEm
kGZKDqu1/qeA99v4zRr19p/F5wRmtgjeStS7AC53TlaCTmAF/QuqtkNqWpsEP4aJ
U9Qe4bKB7H5mgiKxOSa8tMRwQd3d2MvNDDon7oDBYTlhDDdllFceIFBEKPV/qgQG
ttSVCiubd23juKEsC8pdU8Gc6udrjmyjEP/jtWmtjoaPxcixedaxRTx1IKgB/VW5
6r/v5grR9uT/vfgaTGmh4Epo3YgI34GJZjqakH1799Y3LnNPMtia6R+nQ6naYowc
sgrYa+tMZp4hTsVYUR93XfPx7fQNYtSQIucs6YNfdtxk1L4IBIxwmKOVX8PctoBn
l4JtntNav3K4hQT700QsY4XxdSQZajQTZMVJ2E8qgpCFF869UxfW9NqtT8mT6VUj
ynxvcSEMfirdz19LtzU7X3QFBiKTnyBawiQwu1qw0nZ1oN30WAlVjreLKnHPKYVj
05MWP+oxWSnzvBJ9d1/L70gv5kwq+k/nbj3CIx6k5gDqIhG1RbHPMmDRZSyZoadT
dIu6TyU90LB1Xu2tNAoxi4yqAbC/HOLNbUYzFWvw2imFCXeoBZlno4mX+Vwk3gIS
zDJCuv4koRBthNLlfYFwjbVgtQV8Ym3wlU7WZZ0bF2L+1DjkpLA3l8/HbDv23ktx
vBOlcFJDyss0wwGH+plvta2IhfOTfWkPn9ev2jLZYG/NScLtJghlHLTg8Cpegy0w
SxHZ3HMex4yABEj54yLsM26MqJrwUbqvvEEs+QW4veI2jkC7mLPKwCgEa2un2Rrv
mdZnw36LiO/AlonZB//KTrjWhFDBfQweNuV4byyzMGg6UfkYs0BZVnvXoB/pIECF
74W1MItSsoRZc8n8z8gCfXs8xB5UT4TXuh8UtI5wTAyYMKbrYJDhFYxMnCIPUdeY
mXp6JRAqT8Wa5Y3bn6isl6u8H8sahKipfhwmbB5bg2br1+FlqkOZtjmngj6rTeAe
TMurRm99m65EutxECXzU7aSeUACmu3FhKv7osdwgmdapvrUDRNX83pkA/e3V8DOF
qkGXkgr+era6f+rkgK/RwpRD8YrMY9NsvfsO1oZ/QH7IdfWXHm0tnlNnQpQEbIuh
8qSs5eCSTWcDheW3bOijs7V0YUBBF9LmJ5N4O9l96ryLlHXauHXsQ/0y2p+LP6Vv
4ipp7dOWf7VEgNK2bzopRUjQUE6JilOBM2C4x9Wxs/xx/egW89Krv6ufOKHuYOHr
xoHKGklg2AaiWvNHkO0AzMHYWDfhS9PhwAOtle3tgg4Rn9SgIJsNJBykvlgj6Iz1
hMP5K9NDf1+RG07w6rykcjouPikXdSAB6a5pU3rFbDjAxkM30S5JCaWGfQl7wftV
gquV9zG5PAq1QVaqodJnZHM2TJ71/GTeuo8tKlaLgIdUfzOi2KkjkhJBkC2VBsbX
590PW9sgt54N0JvAAQ1kpnJGIAKWwhwzjF0WQopvvP2en/LbLpCQACQFjPVtKto1
U4crMRwx8RZJF4k81fTnzX2UODi4mfv15/aFU0GwLEEwKFnFHGbM414GnijMmuaX
rZZhWONcRiOkN2wR1Xp5MjJN/TDRQNlJfnfq+0KFyCmf7FaQ7GTtaq/qJwOMAUYn
yxGSFbFwbwKgULGBO5CPSJ/4fblDJCT5ZF9H6dnLQJUI5+OMkgL2cpvVBgDzsELR
tx21oUq5z9sMdsut3wSIi2hF/HshQGdK2VWmLKX/hUWzXAXQonH3Vu4BARSDptOb
4qLqUk7iKfdjGu+len31QVEzYKnNgj7M1xUnHyWk3ePhQXBvV4Hp+VOLiXsPon3K
Tt3VHPmOoP5K1UqY7Eqa4gTKKM2BRFUVPxaUVwI91CZDhnHvtG7yzFuPS5Zgi/qb
4j+OpTF6tiOgHirnhLWSc5LIuXZPjsW2k8L9E3NdYiT92RBgrSwQkwnYCYRIgugJ
h5+XWUJJkI4h0fSXkQFNSNyZvnsycSv0lukhanxf6F69RDGfh/5NTR6DRZjuq0ll
cQUVZZ9jqS/fF8XxZighEH7HwCevcDNclYnWijWa/hTEfiE3TP9j7ZqGdcG6K5sk
QFLwo+sUPAcT80iUE0slPjX7rkoqfuYL9RkL8m4pDmDMNh0PfZk9Hu3kfoNO7WyU
1Vb6Th5AyxqeuWDHzkK8T1odBDkwA8OU/5z6eNWnyuXC+ToXPPF7jyQCJCb2ywSQ
2vGkdr3rLCJN30d7SdIFWWK9CtFXFxwKiEt9ftV0/r1MMsSdMhMTJdsvZOMaMAY/
588aEzCLaKKhZsCfIr2a0CCWFYH6HjEqSDSreQV/5khlcu2CkUg/p9/UE2crMpLh
heR1UUP24Z1Ebz3/7jDp1u7KN++XDc4zSKfRcAoTJEpaZRkMraEWGBDF6X0n57LA
NqhU2YI2U7DVxkhFo+NJLvVhq3KtxrQSzqhbAp5DshnQJdcht8LqKQ/MVZfO8pz/
JTiZn96TcENE8aR2RQCP/ACPQ3ebkPz1Nelu+U4Y779XDQMtDOmULiFm78c9sF5C
WkJVJXm7+ooNBza3y4JM5a4/TeP5UoCYyqjad+11xZTllvUnqVAE79YJ4C0jSU6m
t63rqOG+3qgc6O91R7nJ0EeO+DgvJf9tf6bN/RFhu/Yi7ADu06Py/Ffkfvz0s3BL
WkEUgmVqEcS8fhAHoz5kLJWroPtGcSlu7fJ4A5R+a9R0bjNkFzHzyl/9ImPelsy2
L0i70wKeIxBlD42RDovv/h9K1CeY3IEa7ZFYi9TGarqNaRsJZLTbgTHAXaWEuncn
RmN5AoPNZ84AUj3f1yB9GRvXb4dq/Zt3K5rKtNgwrzyLRPkLORVlIYMpXhA/3WFF
8aVAfFJqcGYqrnG1diCTL1/2NCqZcPWObbCr8l0tW0ZCGjWogI/aWkCOWPnGUzTb
n6kMIzuWDBxIZ06jg+w8CGlI40kBEV3zdQfKAVdpZsB1BY87xVwdmujiFS0IhT2N
lmNMEYC8TesQTWW4mBbMaSjEqq0zsdcXjzUc3yikqPobHml9J2tLnJnovkCy7RSZ
Nd4gz1xom9u32R6kuI0vjjSGPf0nfBPc4eT+DLR9ehlPO88RREcrVKW+gSWaH0YB
Vu5R65/i4uJpaZwoocqgu8pUtPyCgV3pkMEaWBGIzzwdkKmuH1USF8TIbf7CuxpB
F2STzuEAGdqR8P6iY/JiaNYHXqcOV9E/c9sCNpA1BmhGmEpHTSwGno939re5RaOT
bT+WpfntBslOCzQmhAL7IDK2fsV38tzZwQ6pksgaP5zk9kD/j9s0m4PKrzE0HsuI
DHZJkiDttbg0mz+SGbtoxcfp7fq/PGvS4FLcAIFO+0ATi0stpa/VaTfvSbTvVpas
WjKD8VQUG1i8aKgMjuMnWuBoML0gNCRz/lCahHBIGzs4ncKZjcIo7jRK1CHswCq+
h/e9Nlqi8241qVLY1kJzPmLVEP9GlOj5saii5V7Xt8lI9O7PyUoRNqsFAd+xovjw
camXEIffpLpy5BpntCbf9v+4q3qmC+Shy/kTm8EaLCWqEEznb0mWDVtRXCDCQBKF
y5L6yRmHlexP3OfUxnW3caFauAikMXg5V5zWjQwbVtxpgR3veCJyOv75I3Mu/7DR
rb0uy7jloYtUQHL6BDy8cdkgBlFpQGhpcFbkeuaFgoYOsU59YBuk1ZwtLT1LQNGa
7E3AMe8coDU1Zl1Z6T8h0dVFidQe5XjrR/GfWEh5KEEOYMoqTb0QOwLnYjqJbeng
nBpYRQqW50yRSoCnLvlr3/L4OHr27Q/71OvftJVmOP9e32fPAWHpVC6jXpY8GGKr
FeQ5xdKJTu/8TXQUzDCJFLkwtGPTnWp2nnYCX6oc9CmylaFR03t0mMhCJ1yLC99Z
6QCeC5QfK1ynDhEzJFaYsxrtm0rkj4cWCz/UeNsnGPw8p9hJNAuIhnIFCKMAfzXM
8/lvNuYH+HW65EkDHm2M9v0XjrefEWvKSzDmBXH8bXh/51R5IdGlZmnlrwfi6Yqi
+3zJZcQ6E8dD1aVIywrFJDzvnpxtztNJM2DGOS6NPHtZ55rIKB/Q9IR/92hGdAbW
DPSrfMOJziJ6G5ss3vZtZzkmuMY5LPqT8e38bNkQY19DpK43EMXrh8dVV0/km06Z
qH9TnJ54Ve/OamenkPzSC9u6fenrpfjmcY034bGzzeiEdAXOZRCyb5o+SoVwCJ9f
dCe9rddIkNuXRZE5YAKLYx8EDqoaDVdMxTgk6UTk3BALFKlmPYw+aO67BLL18I9E
XMU3FpSYV20uy249rYrv9IaRiK0Pab2XYtzwR9PX5OlTlkNzGRqzuH1tqmRqQlM+
`protect end_protected