`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 2016 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
2mA4eiZXfChkavClTs5gUfMTIppeCn3MkfhSb9uaDxxmeutuqUHOwzOE/m4UCuCK
1JxBCjGAN/kQpU+4fXCXHV5XstLL3f0KAXWN2uJZf0xmHiRWBHMJoGmmSqY6zTpl
l02bPeiMkU44ePYiR2usi7/oVztYuSQlYi0gDfU76JEiEEuzdEiHPATIqWdllLkY
p8ptt77D7P5U0aPJO4jWvNBka1YSDSrq5jKfzkBLe/XyGQeVm61vo3U3s61xAnuj
mFhXwF1pM59jnXCxoEo5Hs4ODWdzysf07MYHgsbvvR0kbz8tVSw9tZZiaGy0D5vm
Z/Yy7RYpZIJVKzTWQfn2vspx+3r5du9LbivJasWSH/0QBxZGtuvstIqdK+uzmUbC
Z8EWJophB8qEKgvpmaYVSipPb4ioyMImMLJ/Nl+CCHv3U4xl7mO0lPuAQxbOBOIC
M7IBeT217lL0PIt+9iaATpZvEaTZel7EFDa2RxtR9liirtDgConnIbUJ5RKbmH9O
uMFDPQBZhdxcJ1OOiQUeV86aDf2uopQFBBmVl2dykfW2LufX9fgXCVXkJnzen/Yf
8P0BlTY9inrLGGg53RHy2sujgNwsiKk+2XrsY7wKe9hJnFUngTPmOBNWuZki+zHY
AEz28aW5kiUAfRLs1rf7Z+R83YA8UkNQ1Acq8UPSkp8fwY+T4TXEo1/OontIVJlX
SWq8bNWMNWhNEske0BECIVrMD0RD3U9SvX+GFIhuouXsKBN7ATssQpxjANXD0epM
uKNnUCbCD/CSfkCmicCNvolMafk7XuMMjK92NJDMxh7Ek9ejsWXxjW0BIYHfVawE
UenZKxk36BwEVFE5DatDDt/lFkyL0E8KUDwEw048u5qY9J4H5H8CTPyy1xkwfvTI
WbI9gDWJmF5xyTKhtuv5O2Tceqg0p4yaxfsyivTXRCqXc0zWMEyjdgzyAwkqlTed
Vf2F+wOT/Jgj/onCOoYeusCR1/I19H7Mo5h5hJ7TmA63VKFRa/rDwlbEzCvdqojx
jojkEM8DOds65MIysga68VuQVKJA3dA21IarwpNRga2xJVMERL9vtzOHqTG8M8fU
YM25XnxGI5KFxeER1FdQAkT09nrGjgznzt5nSVKsOTD9PTE6oyyEXEazYA1LedTv
Kf4NbEu3fw1uCDbg0nnth/+X3imjaBKz4tl8x3rXJxR0w7IX0KztSSibZh5kooiD
y69oR6yP/WtikYcKzlzrmh3HVr9miG077NKBGQ4nxDf89iUbLylxoVSA8V4lPUM3
/xLHA0sxsvKURFf97GnXaoejnF8fmQLnJw/JOcacEqLIe5Twq93TpaqHEP7S133T
kuuA5zncfqC6BND2wX3K8WCIzoQxEhGE0ts+kYsbkbvmiEokekWT7VgQmbkvTuPm
nEAKVF/Y+VpPlubUjgzO8qvjz6TuOcoWRehJc5rKKlvQGknXfVhnOMVEGNCxunL7
g6rcFPFCEAGnJUc/+w62AnDUHCJBAlJ1+66LoMpRG9l+mRb2zOLcq1CW99nSoUm5
lPkA5OHvQuCvpb9MG2/y9jIgIHEu4gDY53xTp/VwYFuP6ZAb6P8c6cSqbArqyHJb
Gscvhj4wGmc7HOKXIoC8KfO0UzbvoOjYJyADHwoIeklbqg3RTAoxZ6W5Pdcmuv1E
xNpPwzTiN19vT1VrIrlrX2GTLg11LDzNBJ9SCIjqORH1fMXA5UCOLlUXmPSrMQPF
kKfrA01Uy/FaopGKU6ZPTGssa3uLw3rjRG/ZZ8ayLtSn+UxVDRMvOBQGh5EnYnN/
pqS7A3nx1lEUvqfv1qVgIJRMI2VP2aS7UD7173Za7SeO6M8Tq81iQb6fFmv+y/21
8IIAf+5tU87EtbAWHhnXylbUCKITasKqikqNmOznS0tMlLngTo8mcuojBwICUf2m
XS1vIsyPxQ3KLeX/Gy7Mpy3uE7aceoi1BUmD4XQd68IByU37/10RrI0ygaj5yVoS
MWgjiKAQQTxIDaqyWRsvmBIl05aMkLWcQ0b2TkR5yy84LyegzDy69svGgm7wRXgJ
nsesBUf1wlAr10Ok2iCtH5998E/tqZdv7IchfAwPwcoz3kYGkNRWirXHsqT+HPdZ
gaYYElhGNKywLr1sXetuJx7NyTbMVb1AToP+maUf8bE+NReNYKrs3e05EhzG3mpk
BfEFuyDCG9BCTnb+1OUe4UTDvMNA/nFThbj/C5r1HVk58up5e8qFoDRVoqpsODxL
dkhD+C6doJfgTMcq/CUVW4r7RuvZJtXyZgDXiLNWjJQsrpIKYuz08ZVm2Jpm46fB
l8HEqUh4t1dkZlgCgJMj7JphqOpweQkO3Oiw+g1LC7z2LQcPVEExtYMKiy2J4YFi
rUUdZy/SQq8bMWb2VsfEQ2E5QIg7VOWCtGhTw3mgfiDZgONO849Faqg28jrlqu8s
tX7tqnptKbuAAhjXq7Luh4IwKDlvRd0YJRGOKagtFrGgIDNcKULJjkNanHIS89VY
79VOZXXHwlFaFb88JAVoojjsoHwDSlx2njrBe7YbFvxvnAnqrUGTEGDhYTWdp/L2
`protect end_protected