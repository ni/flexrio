`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 45040 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
3JbtNiAekMoRUw6FSbjvdFp5fj9nTitkIod40fna/DyGd0htAO1LA1G3JeUaAPso
Y4x2ZuOvkgJVjVHbmJuyUV7tdEA86bXloR0FAJKsqJxVcLCEjoczqkIwV/gU32oy
XqWtwdqDBl/SGpOzlDnmM/bsBr4/wSVEtNrolJs7ut9ZcfwwPGypbAvC1dd4L1EQ
rbKHWNmfyTx/pJJdZVpCdwAK1GqI5lCC8KgcMEdl7N6pZ7HtG5DrhES+os8tXunt
fJ5ygYpqk9UsBN4YRlwQvA7Qn0xxhg7iU+FmSSNIRh8pr6hYIntxWZ9+rL35Fj9f
6nwVOdOD5wGkU+LYnyKG5uDtsjRK2QCiIaiIcxLHKZiUnPYT4/HX9aZJyXFdgBaH
AoZkbL5RY2dvZt27SjHnLw7eAITFzTDEYzz5sh9cSu0icBEiikpdUGdNGtBOMqup
n71Y6S1D7cAeiHZh/wRnVrUCu74eWFQMIJ7Q/hDSn51/GPjj9I2mbaIn2uFTkL+9
2veVUSAc/lgPeqQri+ZIxhkIuNwdOSPdWh344vDfcRb2LAV3EfgXas+wotjwyaUi
3Ad4cCfXyhPlaoVbIMiAE4Tg6Jw/3ux97YpieqhX1ejVZ8iGsWAObZnT/WRbbkqP
7wsaeE4DElok6dscPePxNZQ6j+RCoug3KUrZn/SLHGCvE8zGH0VoPMQ/ng724Vq7
gA4IuoTtmHHle+86PoPFUK229xCh7Wf8WcCm0t9fqpxCBsVfW3MQeKXXmef3WBcO
mkq63fPCwnYCG7jAbY7L/6ycAFVBU2qclQQQV3/JYQt9jem/tmEA/tJPI1QXMWPA
aNgGqmmGTRLFyo5ZLPzl0mhet90sgPknHt0ugFERGwsdk9iTgUGlD7Zk7dXO7lSv
LI1VDbQ0JB4QoNYNRRDwOcU88dQ5M+zHffuQFh9bnORSv+gWzVf7RHzvXprGAcKk
Q4s8N2iHr+4QYxKDPrewo8Q0SlwygBF0E2TnI0GjVuMWloLhAk0nTy3yJGx7Ia9I
SZhnjezDYeawjvqjYuVZBUQ8OPFMMmZ3EMUK/gbul75q5/EXqgBB9pMjqYlf/kQE
C7p8/3Jzd6bWBaVs7KRZkotiduLacLb5roNHzcf8ZdPeftmZ/W10pVYs/Xv6HtLp
bNNu0d8S+9/cFzdd65Wx+DPPeQmm9nfJmoduevMlBbsi4xTufqiVkm5sT4yjOsHy
GQcFk4j0dYrrgA5xe4vjxfkgMV6vpbZ4iteomd8gdhYc7YkVOH/epwDm9jlc+p52
UOMVnoWngcvIp7zguXCROf6Lh1LXu5d4Ba6xXID/iZy6X4jgqitQyO62SZQAs6e+
DIPjlBwpqEFIN1i20ZL1eTT8lvP1U9NFvNci4Ppv1kwalRBUw+tQH9vl3MAzBw1N
DHAt5o4zPCf1lI3E7q1pQId0uEb8aV6zo4Je9o25mv/74zz4jyexIykSZ98APB3x
aZNBg3PcpcQRHiPMurj0DXqSS/6xNBqmiYeeUIgF22EPOYt+YCdvJcq8W/Du+++E
6twpnhD94H2SDUEzSoKMnK6qwsZQs2I9tIc1FJH0Wj0wu3NSix9FFaAHieABXp1t
b/xzq3B9Gifw7HAQMjiWi7QPr+uC/jKRI8GEc86ymSloyTungssUwGjdQvVCGxqx
X3RnlwwWxo14OY1VGuncnl+mAorp0HWIdM/BiFAl9p2TRmEpVT+wlLTPtB6G0NJC
v+m8/J+tt1mdIsYGJPdflRLt6wTQDiCbHX6JO+P6eU8YL92ezisE8V7eYY9zzNpX
kBYsuPrKx022TrRgR01hJQxfU7I1cvK7OmGXOiiscidWsIeqlfBpzPwk4LgXrcb8
90bWlhgvCwDg1ieVBYwqBXLCNYRUgMTjPbziyZenz35HTe3OSnl1CecxkOHZOmTz
YxJ7Z6TjvTmM1ZlWH6XxBwWq8DjfM0Wj59d9OJwpVvdeq9OSXYV47tTx1BHxpdNs
ATwxC0PSqO0VFuR9OR13sYUiRDEGwxqo7fCIrh8suSjksgxwcpePzhYbdhk1I5Bw
B+yUq+ytQBlWsraP/frj4GWEdSC4dJ+23klMtjn322Oo1BQ+MB4VOVeCwpK4um0v
BtytnQCubzmfVC4PiDhErHOdtuMrTS/uKXnD3T+uoeZCA20Zwg2z4XHA7QmpnVdS
fbtzS9LomvG79QaH612D5goi9rm/YW+BlnTVxalprGqWzBQ4ycPK/v9p/n4M3+Xr
OcgOCztmiMfYEJia+m4hlfRUkjN/26JVFm32z3Z/bo5/nBKLv0hdhFkrtlAcn4fm
u3odRercR+DadB4FEBIJgofrUXAgcGDQ22Iqkohd7mvnE6tlKm7wA5Olc3Ifn4aM
BxgaQ6GxSqWPC2NUE6yrR4IhNRPoL+fdDRS+mI1aXXI2yIBMCEWnW0mljWz54+eJ
6KST/ngprlUYDcVWtkGLIDpn/HH79C4xAr/np1ocmVxTYFLFZrNDN2ywwRS1O7sg
+gk17HQPAll9U699q8L+BiKX4Q+MmP4e1yS1i6RyyfHiBcHVvAl8rUT5ooNxjSV2
37DBw8tOI3pNdiaEUxgMpsZ+7oictnC9kCbzxznyAxJ7m6Qg4hZskDti5Ap/pFGU
syFIKAh7XxUh020K0zRia2pAk/0P48i6tuqqt2hm0CQmOG+KEBoEpgpQA4aCF/sk
s7mFt5GLssQyx4rExsKm9WBhCFu977bHcXHggoxSouS8C2GZzAEVEFyCfhRUfzR7
GJhVPzXdNHChWKZ+rAMpSQfL47rRZ7uYc/CSgCIAe+tk+DD/vsj7UQdk7mprbL84
wBPXLWyBdblXmJ6xOf5YddyBj7fLjC2f4l3hebe0kN6DjkvRjMUx8TxTnTzL4kJu
3t4LuquOuykEinwPmQn/eMgzuuVgRGApmamOXqpJ+Ooadfz2yYSQlVyXf8JSCqGG
YJsseB+dU8Lgu9+Hh8hCExkNgRvDWiIbWq0QovvcNz4d+njdnQGeMQ6c5wxTUZwm
dW6D/BeRkSrCtziJrd6aEKFD9rnOQYDWveOZexzE5EEU7S1keynnajKYszeUvera
XCIT9FUNQsBkMW2gv2H9w9coyH+b0ylmWxVo2T/RSw8mWmpmr46Qo8C9uoThWORD
AWo7vPWXBewtVxA8x9hZ7nptPkWWPYLskT7dsT+e7g9053ZZ3l5ovpATWsD4eB5R
IgA5zfGmIt7Nj7taqUDbffEjskOWxutEj/G49bVduSU9pZLZnH8/PD3q4qInbWQK
Hqn/n9tMoTa/s78tAMLuCHae6mSSBNi0XZSVA8FAACY6gq0f0Bpt+GlpozVbQS6B
BCoZI5LcFuHfDk/7De4dcJfKUZqaT4kSxCRNJtuBBYZ4OMdODXoBcoFtOrKl/r73
Nt0YFK308LuF/g6/eDLONXMoqVWA2MssnvlYbRltyPsYb3/dBpmEee3XlcWOzwr6
VloY/xNeFsUMQrNDbkNl08Qhl6XQXoBslGVE5zrXA2j6FkYRn1yO+EgOh3UB2rUl
ULuV8/hdeOVOc8o+pJ2vjuCcnVcc0LaQT/C7v6U6TxIimxDzsMTN29IkPVkTnxWT
pg7QRNG53PDsKJv8ph97yvjUTn3CTpjzBeksKE9jvt2Vs2n0te4r0ivvWXohWmY6
MyN/JlPelC7YaSv/WeYd1aEGKLArWheGGyAyVxTXpmaKcIB4o5rD84crGQgMNAzv
DO1EQvBEst4ukhlTEamu/InyyZ58+ga7uuEs1ET0S51+qUTFdo4EQ0zZk53lebx2
d1drk6reHPVQueb7R7yB+JqDfYWCWBN1agQUU9wr2vG4c5vFkWR0s/xGnJsAjKIl
yJIXqf4eR0zPDkviojyp5TT4TvXV7HoH1R3b9qJ/jxS5KRsqGg+2LbcMBMDNwss5
liopplE/Zu3neQ0M6tw89Wd/RcppWa9ZTaW0tPrQzuiJr8Bu8flVCXklO8Vb0U+W
KVdTyZL/Qxvca0dqaH6CS+YEBzPruBrY2qzL/rA9rT/pvNfSS8x1s5YKDukTh5O/
0fny9NKR1F3Nxe1EINo78GemPu6+E8+TEiGUVNbEM4xqxitDae60OKTF2nDd6lKO
UKkYkZ5XKI6KNS+dyhHqqeI94z8Ff2CbiCttd82hW2J2EK04rcbCuz3Yk5kXKsez
ZDizRf7AQwpAksZWPSKdNlaopQYIexBb1fVfD1eQcFFFgDeWHF5sLaWvyh0Je6aq
KkxJ312jDC8VWQGytMYTNSwH1Tt3WewO7oLg+w1tsR4tLnr5ixMhGwZMaRecPQ2O
Bj2c31TXP5AdwN9dNjYHgmnVNc86xCO8m6mzEtpRl97vyX7iud7diIWPKHT97vIG
anG4fjF0JUGzly0fl1DWoKjS7j3dIU8CN1ktOYpn72fHx+0Rb2zgEbo25pIItD80
dD3sPuv2vZ860MSikOfWdWiemvAOXJgBr9AutSmCe5zQhnUJq7FGupS2lJP1Hyd9
Q1Z88BDqMvNvU9vTGVX80VJAc+6x7zFWpcleybZT2algDjIxhI6rxowKyFEkUIf8
OQBfiwa+o0HQJlXiUSNwd+v8jilH17D5P6tqDZt/+QeGywJvrFwLh0CR67AedyNs
RQ2TnGJX4+NZDdWqFrnnx6LHzxGCW5+7zluFphSUmviQW0KsI4iS+0Ne2DfUEKs1
gdpM2s/v1porN03AvHQXmh9uCuuMuN5En581XH3oQcOJAKFhMxffdWnm7Z9sFFv2
AW97vJScKq8c6bhHD+e4Ef8+RQGb0OJzleJXkYBsi+7j3EVGHApRDPSrh3VZP6rE
NG4DOg9rzoucF0pFuhg3yYmD50YcYlWvPyxpETNGctW5A7LpGdOb77mJYol9RXH8
tBANOuJBuUzIYWN8u874pGCVBAdVuRIBlTcmVfEMXHrzdsDCNiMUbJZd4Mj39doj
MZqlaTOynIg7INXZRSNm3b8xiBGphHuhNGj6295tBZ3ZLkD7GGJOPLieB2BuY58t
sxICG3k+k/s2Hpf7VI4Ps2RyDLgXf2cDS1ZkgQIgHY8hYHdGAnxAqkSPGfdnOb/a
WGimc1VCajPo1lCJF0cgeqIJWW6vSckx6Y5s3UwHW7QUCscQ9huMd7Fm2tAw9Hq7
yi1rDHIx2n644H+whs90oLBUElMxrAsfDsHIfwKnApPgvdD6niBedjBE9M8q2Q+x
Rf2bqTdlZzTnAdSPrcQIX09TXZIJnyieA6x2kWGzsVoq3vPp5l/hTnQNbFr30/AK
9il8jY9zomQuXf99duI+vHAuPaAWC9YENUqYFObHEePPmeaaYq5YOaRlXvYw7rhY
e5y3ilWYf4Kg9JBP2qqjG25hjZ7pSwt99P7fIAAWk2OmzE+Pkrg/tp29j/8AnJCF
sxXT6Vxc63owMqCNk04kt+zNiWnV8YmedU2KMsqH1cr1ylHsd1yFWoVLSfMRYk6M
5hxEoFGzpm3QDrVpNquHLfCqVy+uFqVq+Y4QPzbRGkYwUdZjb+0wGarvLlJpQs0F
DE6AioJILSWL6jRJwYc6cjeRSM8ooh9/GrMt217Jn2NelE9mnrSGebz/z6plpKbt
e+uJnelOAnBw56ps868GbTfpsi/o9Rz9LnX45OTdpMIuWYvpSmuqPVNd0rMSwuoW
s5K+5GT/4wmSNA+jZ/SBCbjuR5Z7V93IqMOrJ20LAGQ4zK4YPejIEOK3UU4+03kJ
P+i7kn9jw7waIDvsfVoJlolKxILaEZINWZPaxme6xwTcBpy7PyUF2hiY+5cMTWBY
olY4sM3evp/lIMpFoTfO+fH3mGeEzWqbXlSHvBwWMGK1GyZZu0qR6xiNrCQIlMmi
G4eHqxPjr5EEtRyojbbSEy6nbUI+6B50/eOhrfGoWsmdlJuyl/bIurPkfVmLukLz
N29AFoMyjpjGIsYy04fE5IvD0eb8xKAX7KLirxtG238JrNDUktT2v1j50/Y5rDc0
0yUtOANPF2JR0JIGThoXjI8gRs2xKjfVqi11kdDrU8n8pa3DZkhv3DYPm88hY7tK
RYgyz5FKgquNqj41nqMXJOWtqHDNvQnDqsQ0cVIhaf8DWKUFrCgfSVBCQKVOV51H
bP3DkaFrjDlY1V9IlitbzqwcWxcRURu3Z/UcNOOyYRMhd3vP8X+I7eScJXhQ2Zoi
qY6IAiAniAviuZ8GaT/8yrfb/P2U2suFNvCnofMAXi9FWRucyHERBUfEWFjrFvvC
I3sNZcMOmdBycYLpp/2DCKsmGoHtFen8o7SiahAxcO1eZMil2dWPw95zKOG2OFi8
HgrFwlLKAWS/QtkQc48OC+fxXO8omQDLxmcjSvmQn3gQBtoe81yRXemaMRurzMmK
k88SpfwvFRo8r0zIeAKWRG7zg+MmhwnUeFpwmk+mPC0Hhu9fs0wwdHIFYP1iVLjJ
58BNzopcZE2PYFYq/qnbv8Fz5YcCHIwaidtvF/r6R/91GcTUho8EZhcfTLnul3/h
K51RzguarK8MBYsdHTujodq3SXx1oF2d11Rac1zP/KNQd/kFTRm6ICVwUdF7w1Qm
ty5YycjnN84+cE+zqBplJmCHxqzDJpH9SKdV0+bDGJ5fSgUGdKaH5UjIpPbF8C+3
ruQfzXDalGnmLDNx7ZOPihm9MY8rUMDVBH68lS0qRoce5mx4+cqmdZkK+d2ttGsc
4Cuz/20PGbpoqn5w29d3XcT/UvZnfpZEHKHUEpAUwtxXH2yihEQgObrafJdA4pkp
7i2Lyb/rhnd/QsS9R2Ux21PIP6qfDf9r+OCEDN+Cc1p1JxipnN4AIcF+Bx9EL3PW
tRcdY1nrWQun0XZ7yqcKLxta0ro663XwiPBZOURlHyboyPQTI+e8RKD8BMB/SzeG
k8TxIPx4o96dk2Y9iDJjaXTzinWjjBSC8SUL3Z7SIt9SK4v3crRGhoJeUemdaCEJ
TESD/anJWXj2jvBJBa6VgpVULFo7xzePbe1v3W0A0yPRQebLQIMPuSQIsK0IrOd4
sB4R7z65oN/HMXwrnOJXDHkkK2adMsxpBYqusbTvZX83HDY3sZYvMaNlCXlXbTYY
cD8z05kDTLeAdaF/LaNuvzzenkTPMQJXAoTKLVKIHTxtXW2FkobPuc19iqth4ChB
Rh1rpKtjeAGyNB1Svc5ndZnjasog5UqGN9VaSKORBQTsMJKrZ01+SxDKWmkAP724
RzNMcfm8PyVLyNedfGPAznaRDT/fApi84J0bz5m1uN46efZbROZ12fR94hMKwL3d
1Dv/1UHhNaAs0U0RDoG5KMsJp+Wb6naHx7HcfYb9DQZfFNvaVq2rqwTTA2haJB9D
LeedzAMsoy3aySWeWTGYIIa67F6tjqCvaXeKsLzbTtS2Qb19igLY19clqYQonXhu
J+nhrzIUCZttC4hhwMMI9ODRAwN6I4Kz4YOq+AsqgLjLTSvHAiNj+9s/wzL4bi3K
rDXaohREN3NzXpIk3qkdms6hXwazIpGOjrWrbqeN5OGCH2J8NtE5e/Odr+nh5FYv
UZFCyKN6UBtcdX0wK5Z2k/iucvJchvS13KUW9rECboGb2CvMoVr12syi7cPupDw4
H4GXR8AiyTQOnt/70qgXFblTDyVf+sYv/l7tX3SJpapUvWm0G8CJyaI/oCUVUhdF
P9m7HqghhEJj+hZmLmiojxatnqusR4giUljeux7o6DGrR+9drlsGv+Rs0rAcADFG
vbE/NRRFunPutVNFja0kPUTIdFR+jh0Ha6RRSaa6HQ7eoGOrbkPsZjTLMh3mse3k
Lyf4eTJ4Exn5onNEDBAuECnPMOaeLi6irmE88TM3PWXxC8hlsYzclWpsqzUoGQyh
fYRSQsasgUIf+DvnZ5/AlsJuk9zuYASBzBH+nCNzgEINQ+ZESAYpwembsJEuavP7
lAjcH43uLxPaBP8qxwhNHZ2nyJDZooSZsmFtyZS6kwbfvisV5bXuy+m9aKA6pIjf
YTM/gRKNye5mEfTkZimAM1gIHtc42Gjmc17f8jxes+VcPZxrPZtBzarTB485Ysc5
mQxfNkpEyUmUOtfzKIXYP8uSzLqAuEc2irkElv3MAVJDq7fKw0obML29bqfJstMw
xWtUDFcQnyNHDf7NpyKa2sexgpzBLXJB41dZ0F8T5d2aiiNtvjVppvXUyomXCWRD
U3TOZn2jG162qsGFCR3Nq5X1TN96jcnXCUuBH40FEs58hCLHS3bdaNthSradpcFd
yXB82wLGbf8NFU6UEf89bcqcxZCBXOrYdyHP77/b3FdIgHrRV+7SXLYC9QsyBzlE
/oOch1ar9KgKIOmdxIzv371NRYfxRgctwD2t1y9tvTbIRrNMa7oiyIW368BJmBNW
z01mtr3KDMS65HLJqpK9D3lFLbGbdg85qzZrQPIa1Chk9GjFB4QmSlaFdOaHKlVo
BbAkQvk9gUXraTaDRxyhwXryHrLWvd9n5+Gk56DDw/uSk/cGY8eUdmxb7iUeW3Oy
IWofE8jVo+747M5CjeR9/LqxICt1qGZWhSoKDgbHvyqNpXpy6AYRnqRbH44dHZHl
aTnUhmbvmfpFPYgnea77knWwgV1mfvHC7H3yJEOSDJXNA3hh3bFmJTs0c/2WJ/c/
C7VmtxbMd5mOWomjGzhwvPjWztU3BkKD7amcWrRmJnCcVl8+IVHSUT1QJOvZKbtF
688mQNv1CPjzQcyWnkGAvu3+4gTP85Uwq768BPZaou/RhOOtGVDyCyp7EKSWeuhX
L6gwrya8cezRXz2uNiI4Oq6ibbdRkaRVvuNp5YMJsHkH18TTN9RzLQemVC7zpR6G
pXZ3YPShq0Kwh31LOACdmzcmc+zz0vEuakf0zis4XaumwG/bHkfB9gwkoo5WlgMF
zmHl9yuGEfylbFijFvO+Cxh4iVGmSxcCGp2XMPMkIosY47joknaNH1BMsOtYIvLA
Uf/JScrGP21LIUxUU2+iwT6zznyt8TgvRYxIqqeNOxf/Zyq+MAD6Zyknggak86mu
VC18kDyKxsMp7t0LPoz+5Ej9PTNx55eOAIfmA3//ho+jpilU31EgPZ7spKn/Vwby
rRcl/2tgcs9FJEZlahK7pnlmIcxM742vPfsmvlscyozxaGNtk+HP1+g0T00oR5jh
7MekozJz4VbuPLqAUe2PNYZ2omVeHoIq5wpNMnppYFZWZKtHH8KrudH8CC0OhnnX
fj931hTQ6pkDKD9tXuAHsb8xWlxrKdL5KutfJeeW7oimggHFkG0vlTmg0nAfj6S/
M/r51+bHEjJgilncqbMWGHg3zlLSmeuAyxLnT+nRCchwq43RSCJqReDqmJmgGIT1
v/MbdpkpSLYk9sW+qwYtMjC9v375jvtqNRQsRF3Rfxxj+cGYlH8xBKkfZatGYYks
olqH5NTJ5wuAINkWphQ9KeTvpIw0Z2KtTTWnoN+DOMrqa+KeKDvtzWmLktgS2A2j
i2ldu1pBbiLWyKE0UUfubCmyplDOIrv9iQU3dZyretSwRoWS2HRNkX2qMw8M6DMb
I1NLmFc1oYeQ772DQdJKqAZnEqPuWyiXhfJ3Mt2hkDdDaAejvR9VoXjuto43iswB
SM0yAIXMPmCOQ5BjEf7sEko5n4ge9nuuScprGhHciccP1D+iERHjVu989r+zJncP
+PHfPAPJJwg0LWEmG5jyyEy0TS5y2F0pAOVzheRotpEgq1WtmpP2xLuT5qIf4myR
HKaR2lVoAWJfq+7EkRqIuKDTrIFZwjdYMnjxhSFZpA8b8h0ElR+33pnq5Tsb2dq7
ohTaF3gvFy084WVXnbwDU3+mvqzN/MrSXHQgylu6iGONR0e7WZarPaBEqtuJccA6
VV+dQS193RNSble8/oPV40mbBYWh91KiebVuvphEKEvHjjIX6SFm3vM2Jvzdyu9U
VMuxk7dXjiwse8um4R8X459K5vEVp1HVMLg1jSaC6zwaEk74nuO58tB3mvWlCyxg
974rMdU5OU/Uep9Tsy6d6TJ/iCrej6LZ8uAK1peehGOua77uoUmQiLg1Vfr62UmN
BKqK2bFr+wM1K3RPO1OUQHdEFMydbdVVklTYiAZC27q9z5dBjQYWI6gOakBPB81K
Bct+9UNGgoPrq08DgepmqjQLnSVBuB6I9eJBYdgDign3wB03pNq4LB94MHUlPdC4
j4gF2HMqCptwcbTN3RKatRg1IO6t0y+UnEz9jAo6+d025LjRY4itnb92soX9tvuC
OJHLvOFzHJnfZjYTja9K8m4nEJtc6wqzdMj1bU7Yrp8yUJOYiitV7KEqcZVdVXhI
KQ1pnaCO418r8KvWlyufJwI39ms+7uuwa87GKj6dmjV+naztRKKKxG+AbVCzxDas
ttjBOMtp4aYZqiOaJzeaupsOJe15R0tnub3pGHTECWXn4eSR6ksk/vO71Pp8/bw3
EgedJiogHCrqG524iey9r7onz/phjWdPPks1qtHxQF0VuPB9eSnxwN9SHgCqhUMI
//DN9pWLnJjHDA3NhCf8sR5yJARtJHdBUMDipVf8aQsuBxL+uxcmFZhI6NGOTslq
9XptYS4mRBiVSYefGW+on6vWiEI7kf85o7AsW2cp9XLH0fzMLHzqOAdGsZ5z4T+B
9xGa6WqcNVmmX+9lhVXA1tgT0Bur0ms0nr49e0jg9YfXliIlyGP3GOqH76E8JR4f
IKt6k3lPdmOGii+tcjlGePXJY7kc7xcKK99RbHtHPoS7B2IHCayClLcMp+tsStrf
F73Y93w9fyY+c3v6xa/Chddw1w2GjS1x3oXCTm19E+7zaB2aoFcvSH46PhY30dvT
kOp3VlJj8J64FhrugpKfzlcx8ih9ZPcK/+/vRq0nWA7zCpeV0Poo9MlQzWiUBGeu
JVWUV1FksKesZeSKRNZsj3SxQAe5I/TB3NmC056Li5ZMx/5jXSZOejd6TDYZaUBA
8A/dBMPp0z8DyH9DAw3WMVBArbc0FHLgSMqe8XxXdU5O5FRe7qyceQzXLEOQV+Io
XtctCkyT7L6uTBEstDxHYFBmZLX3QSHkgbU7V7aTCW/Zj5NggeNCdn5TgYB8lfM3
9C93hu6ILjDPwkEbjzOPuU5Qk1HisoFrrPshefL7+7eRZLXrDEEVZsra/9nFIjAI
XUOyEmMFOnFvVupBL/CuZZOEAYtN3jxoE0hytjTOKp0NBK47xrwhLekD4NRSDY7K
3LY+TAfyrQVEa2ox2D8rpYoDsLV7xeYX3QFJ5jevtV8FttN3HT7/7N8xLsWA/PNN
RfPFCuT/Cxfs7nN7qso6D/zARwk9SxjHGh2e1XP06RT3jtzNSmlKZCV5b7EgLit7
CJpXzAqifaFapsUPZrfZ7RUoVzogdF8aqLihxvoF8Xej4Kns4MN0TrDOQ0o4zDAH
eBCS7dI6G5yzz+ljPaL1HBl76+FAdJe9cS1ovCE44yOatj2cT6nvXm6AAfRpx469
yyH2eIePDTkzQuZWHL8rwpKmZZFl0qxlB9HzHIjpT0d3jJ1dVZ0MSFSzXY7Ti8r+
xcwPul/fytAxSP7LaDmELP8gmOTgq93N3fsG6k6C4F0zwOI9/9TQ8rVrNVvGhvCf
TwRu8X5wcAz0dcS2PJGupiAb2Jni2p7hA5f3pdxsmKcawQ5nTj6gYQFTPhgtEXtX
1mTQzBuDOhCtHYps46BclRNdAPLOZM/VhzO8C2LlAqlZ7E+SMUycOdz0uhqpWkug
UKDGPAUhHVEvFce2znh32VC/2QuVHDqWpNx3c62UmRSDn1FlX4Z1YY9yiuEzKgCt
mc8T6ExMzs2Yp4bQqwVIBV+l7QCydEKnUQUnAr91G5Yjn+nb3tWuPAUalqugiKNq
29oguSwnaoUiSHlZE5gbR9G+iSaQO/EgFjMWTihXLpL95MQMZy4IymU2KKnesBdw
OZTbfQ3ipPAS8mw/YltGx3xtZjI9d1VPRXvUI7SAIK5/CH0goGNkzqxpKdTZ1mRm
/d1aLPritQRuEliaTYTr1mC9KSpNVAO+swoa22d0Tj/uLfFPs3yeZXhZFMXbmlkJ
kz3njzZdU38jDKhbof502Kr1kXsPfSE8PmPqrQ16pazt/KNaGa55TSIZLEBtDlKc
YPayMPxoxT5H3o9Y5LuQGwzkRnjKUlsGsi4VgrJqRrUW7I1HjwqCfKh0do+s4St3
/SycVZJ05K6Ri54JIHVdMPhhGkKLOKt+I0B+mjcEplyfr3Q0miDC57NqrL+bnx/B
efdktEIYLsyRWLwAwn+AHvjEVAdzKgTdw93vfy88r2fr/wgGf4A+T6oW19BRTbtj
PVP8F37APg367EA42YtXg5Rq+OjnFvYK5WyoCkro70vTR/WALO4a8SeeEhnn2lKs
NPQemzKLbCqoNCWDwWDn2R0mCyFy9/CkRRQ6alWog/4vnP8WaJBz517585BS0aJD
xHE1fftocS10MvHlzDYb4wGUI8YQo1/4wiX9r5VJDUHzZlzEAUM120jTPcT+sLYE
b6wm/RThxxeXe1reODA4Rtjnd2iaq6O5wxCdiJiBPK+UAF3gqqsDJjuSUky6Ir08
9Vn17+kDTYnNKtnCA3gim3rYltwMVV7x8J0WZqS/L27uXryemsYBU1uGoVHaxdcr
XErLFkgvqJ8QNNAfCNLhgUL5vXxYqA2d6HDiyG5+iWkD+vYDKJqDseCZS8jNR9YW
9wz1E00Yj2LHsW21yKFN9Y5I2GIy/h2nm8Fy7+NUBtpBMbmir3OYiOKlg8KTCjU7
U8dTYSCXRjVWfNlSGik4xdDd6Xyk0zNRjyfFXtGRnB5DrbteYZSE3RFUhLB0HqH9
GWauGsSS9wPBc4e/wxaB2Q5SQIsYrPEaxbAT7wa6lmSBIHThSPf7CgIulnl2kVIT
u3G/m9JT82pNl467+iq+4MOdp8wyWN9C8SFBP0Z1i+e/+KEj1fX/ep7cxoEcJt++
n2s5VTvn+fScuNcMFh5ONAgUOkahpn4QyLS0PjZrDkBRls81F4ot7KUv8VhrR9Vt
L2/VuoyEqtacSbN+JY6Jk9fUOLgwuIV8iv1TD8exfZ1BI6DAnbYpe5BOzvQ9PPpg
HDeKRT4qG0qtAnSjw9PoHqySOpOwGYKLVeWsumIgtg/AzIQS/Od1FPGL9w9uvtgr
4373V6BasOSMGq6yrdvc5Pwq/k1r6OU8ARC5qNpNLUqWS1fpdAFMOFL+PVADfra+
S8WPiPSmXeva9Q/KhCM400dsPowejn/6CdZNfWFLjCcrURoMVqX4MNIlOm2ZYzWb
zSK1wmxMyf1osRW9EVNWKmrD/r9d7Z8+4QNLOTyx2O3wMyNydMva3LEdeHqbCdsa
8AK9+C0xZsEKt0Kq3vsjlXbecRiKpTrsJ2ZMW7PqMJxupmiAJJmGQ2y7rPd0lZZY
IDbFBzqFfEI+DJF1y1Q14v5+9ySY5H8f5GOsg0oIQ+i8KPeSUaiD69NLUou/i89J
hJxuvtofanW0MfGYLI+Ve8UGeY1priO+W0h8RyxwR3oaKGxEAFuvnVKrC2Vys4de
IrVCNgOmcHIWummJbQeA9qdcmQuxTtsjPo/fWvHZeTjeDgtTt2J65S/e48NRM27s
iOCSepVkJYKY9JC2uPpbjTtyjGVxtRcOlI/jNJ75LzM/0MdKayejnV3iNJ5lC0h3
BYIhKFQxv1rXMdhR95fUv1D3lF59rRDn6woJGllL0r3bWTvO/QDSJcRHHvy5QPbq
uPhAL297qn/4M5481bg5w1w0HS7rLibKLF4pjl7YKY/InYg6i4MQX7ckT3pikdmw
WQ3GsUfHfn8JDKQaYIishDPpS2eAVuyX0kCda8pjo/yqo6fF1cBFghAnjh79qhAF
7wuS+pENYTaD22FxWfLcu1/tX6Wa4LVoRJYIu8Tiu0pFv+tqPDknQKMyHdc9B1TM
1bO/49z+g7loXuN3ADYh8jKjA9xTN4TmhfkBKq4illKIx3NxEHyMDwpAWc5LEl4v
4X8tdGPoBXvdDeiFI/8kj2xiKG+fZvLKwNaMe92c6liJqbSf13x/rIMCAlxqDcfv
SO8+ulxXjkHyJjlka+7+dsuYSjusgoCbmNTjpR6Ww1pKs2m/bJSpJHTUJhUn9imr
V9WcUvHSvtUZ4GDpWaJMOedc9jSN7LKgvUYo2dA/qfq1sD6ZM15ivivXha0y/nHN
IS70+J/1IqFhHzkyAsDNc815oivxrr8ZrKqFsHoUJHi8Q5Epo2S9+JknQYCZvqjl
TG7gmXLB0iNphch008O8kELIOcOlevbDaZiCyUVU2nEdIttT7oOLSaHgsPO0/AFq
kImgYdwIc9IQ4YjXL2aQaQOPZLln7fsKHqsH+vnZq5xWXMQI/eIvvncijnPS5glS
7VHQfYK/SHKcf/13GUokn4L7m2DPkJh+fSCcyc1ZfUxbeqQ4eDy02efJwRZQ9P3g
epC20Z06nyvxb2cFnejbrmov8tJwKAMVEf9HTlrARIAmDWSolQ0XS+1Ve3xuiaPD
phUd2COtmN3m1kymeitvjqwRYb60Y+e5l3ckDoCXCa7rFi3EnCXP2IZS1n1dof06
dSx0xxpgaKNgfnK+70Job+oSn1nUriE+OyVLjBy/xv+iuDdgEGW6dW72qEjhPWFU
ls+GrZ6jNb3RxTgdmQ1ps/dcxWf+q0346L0MgliE9pWpQLsk2qMQH8q9IuIkXrsS
DmTdVh2jdMEQ9yRlxDNuXPBPW8LU2sI9ofzvjnArnFPIiYjMY7iWRg2+yVZfkzy9
Zt68P28fOj5PjjeB02jJlkoidY1ak+/7cZ+jZrBwi9A0+BRj7ecf0ccNjn4/gBbr
AL05L9ZFZW6FCPrGUwXRPbzq4dnD1WiLrzpjQ2lKpmT+MsHB6ZmDts1uUF7b49bX
FauCvkCRIGiOIbdig9CBH1yHXcYaVKVT1IvcBPiRp27Vfnu37kZa2oCRKF7lBfsx
26RsYly28R5sCHoXE9Kf2j0H/Vsm2kOwT4pMduEJdUrPLmp1PYmC4O3MBcELuvC7
U5YGGXkB0mQDDqCMjhp447K8p5nGQA+VS5BAe8lmCswxwFzsVDA+sgizyLsUxf30
aCTK7JIA87xB7ycnvhpFiC+7LGf5wFzzv86VGaaGHKLm+Cxw7XLXCod6voFUUjOY
zGW470aX4oOOG0Yba31iS3jZWrWHhunQq6uPwZSdLtxrf9KmcQgHYvsJrZ3U/irm
yZNqw0iF5iD6Kln0PMc/hu/0cXi84dJwBaIz3GqyHiZYl9nCMtaM4LdxuFhDYIUO
kaf9lLYMdJCciCLNGeLxGm+vNNXBoTe8m89SqTOeGGBJKWCV32s4fiYaxjH6pkNz
IzieTVzrMXySuC6vXAgxuq4sNHiPzkQ06TmHF8MWcJ+rbNFmgJfxKEGEkI8Ay5oV
ujjSRHN7EryXi1OENPnuMHMaIJeMFws/g2Bi4PQaBqo1VOFMx64+51n/PmmJUyDZ
rgnh5UMPpqsWBsv/6mYgcMWDO6tNRQdp3I961cuKjuYPeaf8LvSk4/A9NqUHUxYw
v2R+1CbuplZeukSLHeNFSJWbRv8mGk1adPUF2eJK3gb9qNJfkSdRQQlmFU+jkBCH
ldoPeCrotTqdauNmKRkh20uZufdAEOQzbZdrTq7nE1aDulLDfgMvnHvnx8vPNdpU
oDMgmmUKnvWcE47OJQQJYjLzobFYoPiCloZYpAyqlhrUoVQIipIUMERzdo+o5fJw
tG10+mYSdM7i1Mixb8FXtN/iXRgz4mP37ciXD9Vk5eaoegCyx1zwNr9ULTKCe85R
xOIySc0Xs48dcPvNZMC5blSXUwSIRSjxuzMWuiAW2xW9R76kniAO/cJO4CNeMNF5
wU0OSIBQtELC4fbG1PSj+B6s7/62anuqBN/zHSJdkaDX3RoKjlLiLrCnJ/W9Sstx
eehH6b0QhijCtLhpl55zmFzQaVevPHqaQPZaH1PqhIhwyowtvfkS1iG2BVl9AaUe
RoVgdSW8YhvUA2NPB8hQvpjs64AwXu3EVj+Agk86cj/1jBah/hnlVi8uOBAJCvOu
cVN8Aso1e+7RBJ8kKcz07QOAXiFbduMORes3S0YC6C2j7JUdqUOnH+uXv6+qHNf2
Lz4zb1FPA36r4BQ4kv/3dqm6ntRN7OjRblicRo58Yw01cnEXuAVfpWCjLYCZ3CfN
fdcO+2fTKxvRcFw2Yz4Y5oR9SFeb4ffdkmNaClK0RvyAOqoHA5rtWm5WF0LOygHP
+kRKcO9T0AxqWPH6NKZcoBtTQKC6kEEzVD3kWwzjfyI3w5HATGe8NCmn94iP2aiY
1Z03PSzAzaSzKdFbBLNO3VcCFFGHfnFmH4Gq8mA9kPyLVGJ80YyF6DsCegdTcZZd
WxWIT1RQnSzuv0A5eExFoyCGnsw7zjDC1AVP0h0AR8x0IeUY8YOOakzN56p6VgSf
BnPWCn34Zgp+VbsRoqILqEMiF81GELfUQvV7eoxTVGIhB4YhSdnBxXC/mMTw0WEf
Gp8huS2nOXVS8jCwbt/4vhcV7/y7akhn2wfmA9oeMNnQhVoy4rFNoP7sWkjjobVW
cQuh3WaDdO2WbogRRrL8/tjH/KXiWGIvEUl0iba9gw5O6sA3cF1DFVjwrVSoF7r7
zOY3BPpZfg+zQm06vnCuVOm/0wAD1J7Z/AGFcapnEveMnhH71x+b+opdZByMg+7/
dlxdF7SMHhNRZrpn4tBATxyKzpqwAzEe2CeGyW11lyOW8rXTLqk/FoREu2OuqWAo
GBeor+oykyeysFTYiUbKpWCMI/kGOYp+bv49WhhmO1V7/Hnd0d4HiOfi8YdnWlyN
hRC7mRES9ClWpCzFlix923kFIlQF2svTypdge9eCnNGEOIlblDHNESRwnLkVxYGl
1usD9kxxJc+A7Saa7mlwsPRgfyF94TZOQLcDXaK8KrpuPWU4m4jh39MXPEeoki5Y
iP7lBryeSc1oDiyT2lOvy3MT+2OLX9J7HjnegRqwrvtfGy2cXV5GTLPglWRPPI62
qTBViU2Q4MVCc/WoTJ6Ba6gFH2SGFy7KnThTym9CvZc5QI1/vGbS4jtYYRZqJPN1
o+7H42El2Q2mVk1grp35J1ud2US1xATY5y5bVYrRxQVyxbrxA7zz7n1tGuKxWWd/
wueuUU3cXV/xAlFGlDENuG1yAa9j2lqQsxF5FII3yhDc7SPPHOO7UqiPjHZNkYfd
yDsQO4BWhetHaYNCUE8hvfgPHshs04Krzy8vOuwF8yJuknahWbIC8yq86PeQ7ozD
3RGdg5kdAxaDXgC/ArZhKI6p+pyq9y9GfRLecCFU6Z9P3EWyB0ijM2ZzNX/x5d7X
2vRz/LYEk0E/QANDyB7M3C7S9JTIzw8fGnUfkIV86uf+yHHgZT4VjeHMnCM4llbg
6SNp3Ku4POIjwUKtl+f0MxNCDVD5bONnUlEq0/xTcpTQNc/V2RmAC9jx7IYmUvGH
3KdoGtdlLPk8gOnzuruE6H+E4mdgvP7ZbzCwxDBnP2o+JqZsTtYn4tRPFsVjx+gR
VCJn/FpvOyIQJFM6TJpG7gyIvA0HcNkgvB1zInIJTXVbKY+NGLXuYZFzyrNrsr0j
ErDuJxqCC546nAvtEMJnRc228ISOx+jObfRnp/yCQBlWTfzKgZTgopnpSJRXDGzp
gzrY0uTa7A4mTO0EOS6k8nGV3htsh9C5uNUFqXEvgiSbLggQWDlcPK8laT+ATha4
NbdE+GgbjIWFFdJLbwSC5iLmvbA5F8chZK6mgU5m+ikj+hCAODdgX30mVflWKdKF
MdAsL4YCxKwxR67DAZK76e9Cy8aLUqDdxvRhrRCaeczvyyp9W6GAgPMOAyybV/Oe
1YcsTTbisEws9xeswbw3kWjUOVNFKytQov6UrvjwyLMbHLUlymKA1BXCDctthJcc
0MA+o3dFwPM0TUc7MLEauUrqkgMmGdJq6QkYOYl632QL6bz2F2jA/PO5v/TpcJDN
hw1CfaQMv0v+VCaosW4OJ6uZNZ7rRrDyKGv7dpUbyh6GbMAmc1v0DkZZSJsDAoIT
p3jaUlXhH0YzPBOFsrMxPO9p3eZPOIUj16xVtSudkAvRRSj1IEDcWJ/7iBg5vuf6
M2lHOQTjiNOQSoX8ibwr9O8bJCOZbx3YYea1mbHFZamWC1C9p2RhWD/wMtR7g1AG
ii598FTSF0eeEGHRyl70Tp64n1p+jXSidpy9kkRzO2i5YN+Cf5Gy7t+y0j5HSPxP
RyvCNqiwJMEZvCnkL8ElTcBDg2Qz9JCYPjVyD0G1zVs0+7/4GDs2KKbdNQ/axIWI
dJQkEygoJ7vs1a5ENaCWJDfWGNsVCXRbcdOOd24geGFjfQ13IuVFLbF0mMb3Ndqg
Nv44IRECaTW/URZaPQnHmR2dkSOcWHLYP0zeCeID3CHf2ENzzZmImB0Yxs1oH/rx
TaPPJaYVttFD/1uHxl2Ed7AYPVW3wo5IiFhiE3lRQhQnVuLN/ZDujm5cvrjQVFWe
IxKKoA19hDrCDrO7Jj8I1DdpCBdldCKQhK3wcr0cCosDVup0FDCi5uUZNMJEEkPr
58UOzdJxkrEcDpRqmYb/O6ZgXcp5WGhIRCFyFGFpAtFf7sKMpUXdY5MQpCGD1FGo
ckJFchuhVySZeKP+JnX28ToZjKIC980bzTGRX2hkkXqPre2lHk9Ki7kt5KzSZCvA
pufbQhOi6EjFDeppniLk64ET9vsX7240fi0E1lT6lBhFfAsWojEBde+7smKh36JL
1IEZgadoP6ZJ51qPBaklDU2eUZMIckRQ+wrC6h7tB7rRShOUlDBoJUjApIe91LTx
c67cwjcM7+zs9WYjd8iIxPga3IOMX+dzc8TzZIX88IxWasdOEb9Tnv8D6N6rSjck
EU2hqO2K4FYuMDgNNipvLujm6NJe595O4IxaTxuB/hY0nBUyJTLBOMwSKCqkWF0H
KDUdwDACS7oc2SCZfP/tEB4gqsEc6f+ehdoGtsRd8wnYzG/jdlwcIyH/F55/hoI1
eZ0FCa7RU0Ax3Ys+EObSvBJfPnaWeoiaSAAaFqV4iVTEPSPGK10yTTEsolJsTd20
DnWouCgft96NJS2M++omcadSPZLjNbTU7sACJcIw7KeWOo8EfArbZNl8ad1mPXME
r/ONCGoftot4WTbBWvbTF069+8wLQV0aZSPdnFgJHBDAseCmtK0ASZIuNjTMGuyT
NzP0dzI4aQyQg1anw2GPdcU1+u3J+Omm0jUlf2eaAB1ydyLdOM/adHXxQEzUw5E+
vviLnssaxpN+Z2+yFtOlZmN4cxji0enUwv+gkFkpJDDBtB4/IQT2JKynruDoUIMZ
aFRELE+MsU9rRZ6p8TwVEG7b0IsWtXvTwNh5r9oS6vGakdgUTucEE+bFgAYQNt4l
GwTrmxOrUA1p4kHQcS1vPnRaLj9FmZVRDIxLcUkrW4AyHy1zULwr/1z7BJLVqeb+
t/OFfkV7Dx5Lol/vQCIw6coRtO3fkG5IpGv7zOFrA5wkGUhum9Ua9m2on0AktgCR
5P+8r8wPrhAvF+aJIHA2bzro4l/CDC5KBfVvGzV9sT9Ag5jPyTIuijcYDP1JwtSm
WlOigOby3hnMHRFMmpSplT3eHtiJaantdYUvGgDNrlhJ73qrsyeZ8UmQIGcA/mh8
p7mof5glO2CMpX9ep4vy9ubDUbGUSnSSbKzhlz20mr6GNGDtB9L7g7+KQuNDUAZA
I8nCgj8fds2NhK535e+FCp+b+Q8VuiOdjqwxvZYsWw6SSgXnQva39vY6XBdjAhS0
1UTJdbkG3DFzVIZzSa/U8ciXT0DYR2hQgpPPIw7mZ3oF821Uhv4BUG/VB/n9O9xN
ASc4I30Ev/Yh35TDDAH8uXyAd5Wo9nyJMal3fVG+2qxwbOZsMqS/HORubyheetBz
Q6FwrlLAQUpxhRAY3f3Ho4wzKTY3Jj2APxWmmaPvqEpRvuzIiAnd6vq2lZ7Ou4I0
syrQbBztduHXGhHhGFRSJvLaN3o0vup7oBh7kT4XJPXESP0VQPCmc2FmymlXCO7M
lHlkccGpy0dQlN3529YT/hjACMVmoiS+VGHhqgzqcmkiFUHJFia59WeT/mUOx70h
SFAD3oGmxMm7tg+vQMLWP27Sx8Y4D4vfxy0lHVBmPkO/YEixEV5SliSaRwTteHua
JCy/W2GznifBNBetX2b+pFPSWJbVMlQT8+SWAn1rVwJJ4h+0gZ0tVPlXGYdGdnZa
P0k8uwzMDDjV6yPZ3RMtckHyXxWZhGNZ28Ads4Jlwdb7bkNf06pSz0CWDCBq1/Sd
fodOmiNDqD5ogDIcPCBABhQU7pl4OgM97HePU/n9oq2xqJjz0sTg54SlqKIt+CXw
A0VM/YJqYSYn+8ZjPKn3A3lmpV/ytmZNr6YM7yDjFd0/PwDjzA7EiSVBeBolxTyi
ulFPfY/BElaNtw4cKyb/1NsUZwdUNvxQdLL0Iv/H3A8gZ9Szl+E4eg+Fy/vGK0sW
4j8r/uEJypmJpYQq8NlCw5XGQWYUx8a/YkOx1YuYYQbcJR05J/5FLfLG4RPWAFIB
8gzwkHBfAL8eduVz804adATrGK+Yjl9EHzPKsBFVxaF6JJxK00eO/Jbq6Lm7p6tz
EXqiWw+f+muVflvE/F6rFUqZXhbe1Mw/sbBuUYkIIfg4afJb9f886TfoJQbHs6ah
8ErHcTZirBll+v7F3YZHPdu4uzrUNbgkkAf+yCYoQx1bjJTMPzR7KhFbxAKCzBu2
ClkstoS5VRtFec6HgD9S2G934v95EcCkF1Cv+qBBJ8Ezj5fps6Mj8B6RBNA4CVh3
kB1gRFU8ExRD2PUVqKrAUz3rvgxWcKqKjvZYc4db2iHiiG63BXm97KbQoV0EjpZO
QR+d8Qui8ltKDFNnAKShdHDaGxv/dvH8zC4EGxPwPoIi5GRzwyNtNE/FWKBzpbDF
FDvWvSXYCi+vpZk4ngnvY5TMyQjyhBGOp1pFG4fKV8/AHp55ACclSk1YhfEr3CEx
wSal3/enec5+kDolR7oeYXBTJ+6tG8IJLVjM5aQJ84DnhDLvkN5oWyW5sRJNtdwp
Gp1tdZ6V0PXXAywE0SoXYLz6GeX4XR7uJH05hxHohOjRnasxVpYuLEIHcW7JC++r
tADi5fbJhMLcHc35hAaotcbCuolUwfSCy9WRA+mZp03lHvSfRWN35RPOgPAkA8Q4
AOpyCKB2AJE+21gKCh1fEADPrIcRMvtz3zY4y+ep5slH/QYL1atAax0nJPnt/z6d
Ndfg3DZlKzo/Lw8r/DkhOjhfKxtveGPT7Wj3uc7DYkQuFQarWF0nIMdrfK0gzynk
Bao8Zcl/dFjsdlnjqPWLRCX4WHwuwujm2JKlED2bbnnibHJ4e+n92JAecpza0Eb+
u2LtHTo9aQtlV1W8mLBNQNvwjHFWpx4VsMU7Co9stzIOZE+EacudFRFcp5IynFuf
985t7uTOdSjJdQFAuoeCJUgiSxCMQZBEAGbeUYaHnhCDz9NdONEGm7990AirqFIW
Rx2DphjTnuXwPnWQ7VuwIBft10SKp04sTdogpSpPVXTDCqIYufVEalb0bRc+NUvk
sWBrUVS1irKNivVllflMTFphzGrqhoZ03RnSZ8R5QsySH+8dvZ+PH9jUmfuIWzCH
GGxuq4YaZYwBDXWh2gT3jjLHEQjhsARKTKl4tpMAELA6EnWw3K2pQZuAxFAHtc/k
Hfwjv+WxpB/08tfrTL41XdlAMdObOKA11vodIEOiXEaXBMz0cF5mqaAIuHGooSPp
QJ+192RQQ3h/WeK2X2e307nCkANcNg0lTy6JD/zfFqsCiJRy1JhpTuluMXTnuYJS
p8WLJxBRlntViO6+tKrZAC81MKwdgmd1iONU+xtjXzN5m1LDJC5zBsMt7X7JiyUK
oBsCetPN2t8LEC7Ndh6tpBDr6Sn/RROFWJnRvbBD8IePB4Ef089Uh/Gd4ciYQ/jL
SdlHP0mzPv+weYqXjt6otW6BpxBkFQaomMiUr+elZNot5M5uNt3u2NYaKABEEJuy
5oWNRIXoUFi3xjwLgSUx1PjWdm6QYZHVFfBGk8PbIQby2arTtKCmqOefeq7edHwm
ZnuBjnLsHLl39Ie6L6Ya1LzjPXb/7q+bNyNFGpcWiVH/xdx43DtKWJs9wKp5wR05
h0W+lE6W5I2quWcVROpgq20VllqgYyADWV0lFu1RXmUYkOpqx70Mn9xXjjWtIbBA
u7aP/iBn4g8BAVvhUZWyB/KXE5VWDheOjERlgcEA/GadICW65Dlr6cDIWOZo4WH3
k+3zA28NUZMFeLKocD5fVPiLBCUcCyfyyrHaXYb8BoZbJSiafygTSz1/SKZzCnl7
HWV3x6HJxpTTWjFK3xKceqDmP7j+6gYzG+8KxWHWSI3MLLB6XiyZRTTrcCig1M68
nAygFS94j1UuAN8QP92vYUOglYagaCGN8ZcFcMFcuGIV+b7EP7P9iibW7rAtdLjk
SHHIlZFbRvGj2ZucRHA1tk44hHmaDAUUDUhpqLAf7ZytWaWYNrtIxMX1/0Ks0Z01
6l6bco6DI9sqjZOb7gXtqpCFrIonkEHhf0sP1aWLBzYJStWFD7f0Xroy91awFTHa
KPlBU8cjJIeKmmsjkpZrhOd6JCw0hyWgnFRsW261/G2Zup9hOp4T1Szvw1Fcl3wG
anEZfez2VzrXl/4inbO7Yl1SjeidToHUfda4nlyqsVNlvRjEY+HmZlDqNjawWUBp
Vi/Edv4qAbqil79jrphy8BlEGZSSsFmRaohvsx4iy6E6bGiIU1iT+GDDMVAQO6H/
IYRVljHZwKpafp6bRrBMWh0GzWRPYMxm0Ji7KlhwDOCPP9MvjnbXOzrAT5IL9Ad3
MZ+BZudaUUlbPDEZWSiHHszlDB2lJBIJ0FaoYb85+MZMpHUdZZ+tejWL4pmPxlGo
aUh0D1GDxcnFLVT4fLRbgGAjKbXhIH+JJKs4yhZZyIy2/ymio4jl41v7p5sqmIcS
bYb6bKQiz3sv055WZKEdFxQPQRVEYwkpbYOSO72zbTyxrjhOZQBzm2GA1RZB2lOf
hsNPk+eewc42Bk5QdogjRkozwxE+Yz2M+kleo7sWUZhQbrcpp3ODGGjfriVjb8f6
9USE8C1idGvoQoRNuT321yB+8GpZvM5CwOG8v5p4poUB/C7IYUD5MSMqVQhII58V
Wv3ArZe0LcQOL9KQqsRVbK8SGdRztdh3g3hJez89TUXXjn5OhcBjFtIiDQdex9Es
Jsdk0GXLyOnKIvIrlEXDwxNaXST+LtEIsloHPj0S5qTh9jiEGez4SLwxzf8395kD
Bymk1bG3zQLI5kp2FyXr384Ko2CCI2Nl58yRaY2xc9E02ojCqeYFJD22c2lussXZ
Dx6cS+qboYzWdl6P4zw1TPyuBgEWrbq/z11UmVVL4RzS1MJ3rYOmkxln4Qj0RlTV
jo1hlzLcYlqMz1OEUEzQNLi7KpXW/90112s3cZXNTejBWC4gypIREZ47EOWIkiw5
yDqk6XQUDdybJ5APzcUWKi7vuZINH4K8KQEOX3uEfXUdbC3qtoAWlY2WhA8FmVt6
kZLFVoWHU4p4iqrTjDtzRE75nVNjBklcQkqZXHIJUKhGuUjfcqwycXApXNo4fTDP
O/lR5tS2PjROKClW+Afb6rzZKEefua46X44pOgezEiD49TLkDwUHXUzJUZJvmcG0
rIA3NaMuarPO4tH+4etekIzz6E9Unt4fH7BgfGtgmjivCJQZoDkv1gWaeb2OE9qG
2RNexw4h+MBlSJeixNJ0xJxHCTNC+XRcOQtsPuVNDsBegINzGZsiaD1TwzpA0orN
BfgtexWxEQJdE8xB+ZhAZjdQA8i1haMlixRWU6WKXDQ58nJbiCTWD3w4opxISu71
dFAST98cJKTGlVXPW0iCLW5bi6i3RHRtWnmIcz4DH8Ic48789qeBn0RrqSqB22xi
6/Zwy+CrQxft/4MxiFgJmVvR2SgEWow9w1RokoBqHGZFD6cg2Gm4OF/sUFUglpHj
KoiejlXXcRKSKR32KHK3xTk7OSdJUpJrJQuenS5oAeY4n83O5B89TRnVclpzwE3t
MQEbhtHVJsKlfdAWZ7hSWz+f7Wi3fpZbhb83l4c7CG0iaEYScQkFr4KMiD4MM5sW
e2TZqSeSo3itT9GaJ6nxpkv5NMYmJYtyzNalPLjBnK3F47i7wvYIZczhJC83A8hH
gwHiTRv1QgU7q3hh8OzsEj3AeLOEpRGo04vrgnbYyVOqEFGm69D6pUKFib9QW6wZ
Ugtn4Q6ZNiTiintT9imvXKokxsgl1IRKi/JJ/fEfCZ4oV4rAOpYwgd/NcAQbVTJC
wFSHyq7viEVtUSVFOyZO4bdPdX/iTfHXtOWHDGC0GR5+daqeFdElR7nCU1u802VS
EnttrNLJ1YhJC9l7PWLqcs/VbXJzpp/zw++SMrplMrahwL7q9hLKwfg4echzM4tB
QANXs9+GcoW9Eti4Mr0ut+j8K46u4PHRs9FnyHzs05FsfzzMfjrzHOtVsUmRB2mA
Jst8gzMxieMWNjEo8oPEewifJtru5hkRU6INIFiEz7AcvLz46US4Mb15rq9wv+H/
BAbn35GVu54NcTqkBVVqQrZ4NzWL3QrKKco6OXW6daSHtrjCvNVpze/XNS48lIO4
VDQQsYcWTybGpkRG947A+7hHmTC6wg2ns9AFMKpQNoPI2OMCCh9NwEgxjsMbZeSm
cl1X6Mt5OABXZOaxktnEiDj+XaoLj7v5j6T1Uf0EL0GRMdB4zxLSFTII2oq5MwGS
9ts7U8o4SJIuh7b0opAaCXg6XB7Kjh4b8/8/f4Wd3+wFqBLwY0mf9t6pAC1AyCp5
Yu54mNSGahtBJk3aF73ReYpeotWCmfDncQqIfILkvDnP0SC0nJOqrVzTmwKb4/BJ
k6x1ZZEmoBXa+5pitn1M9+KuTGbXKUjs1yElMnh7NGL/lU2ISzrnAUhLg+GgBzdm
NhlfPO6MDTwQhh2yI7dVZ4fP8teHWGa1GQ7gIp8BSt6tDNPeDDjt/tjjqoQXTxZX
Nf/uO7ip8Lrg8yWTKy7/3q5a16EUKfFCjPfrw9PU9j4z4f+a6RUITfuYkfbEtne+
G35o/y2rMvYGdvIAZA2OrrcFaQJFKaWbZzcao7xzrncPNwRM+2H3FuWHlcFYCPGe
xraKRar917zriC8jMozCvqb0z67zwfysHgQENeoeE1vLSGHHXCoGuxcoE3l5gmEX
JFLa5Jws9i/aLDghbG90mjMXBdlA50LYpvA84erwjhdc7y09okj5foNlxA20TXg4
fNF02ufyo/XwbmCKMa0o7WP4voDqOFbYAPDksOODt7jpLDb2SH/cLSu5qaf3919w
I+wcFI0NU150HXxxAhATLavRo1l/0sB34YSDAP3l7eMn3Vb3lw9UKW8gjXSQ4WVt
olO5I5P2Br07nPPqmCy++mzrgpw3jc3AZhCIpdJitrrcdiKd6cXHTHjLtw6iOG75
EQ6tfwY5o9kTc66Jt0BRANo/W6Lnx5bJC7At9HAuoT+wip/nWBJkPu6omc+kwAEn
n16B8ysITI7FcoVf2ME7ldypxPpHEX0fBwkd2LpYI9wxJjZ/uQ5pSeUDku0+k8Iv
ctDI3eprPUCKyc75/SH73hL2t5ibBWNIYX501P/3I+tQNKqvVWtPCVWleDeDozPB
hxl8BgExFSVFRRKg2bMnDm/BdiPBdw9VBwqpn9imwFdhzVeh8hYNIAHOoEBZOLx7
sL0Z6+zuNuO768hdWP3NXEVqz3eECuX3NU2tVKJ4J0p582GG9Bse4rTSIdX12Ht2
LdEqn+eFEsab/5qKRQUdS/yhiBG0J9PW/EghlO/K7VdmFdiY6KyAC2YeRozs5Z/s
PwHw+bVhtYBkdK77ncJeU1X6P65Cg0d/qYb/n707Be/8pPSpMvGi3Fz3AkhAkT3O
ov8j82InWiI4u5R8vA6tAFD+nx8ijF2BwYG/adVb/sPde+UcLBm7xniSLJwSG0fp
bjgN5GbFn9C6KfT8ycYRtx3qHqwHM5JwKIwwbNrvUg4GQNKizhXIbrMuJdyTFrMP
zUg22vlE6kwevE0LPUkgmmSkKaDm0T0b0CTY8UPl/k3aZ+/7zPGCtaHYhQazcdPT
wiDAeTUPO1yV9AMpWaRpCFPwmk+eTG4jz55NiKSHvJKKQ7mn43ph0gCuo1OV84Dz
ImshMjg+Rm6WaaiqiZlcUUGoeoYdjFoqW0JqRpZKMDhEYAT85XkGWunt1Or34+fk
XjLvpLJQV/Te5+BL4WvzZMl4XOpotBG8GdsojsJiBOxqEuF0mxV0Ibr8IYP4g2KE
/OWJeqSXzD2zgjGISURshojrMV0NXDXmVKpKu9rNCEcMFiYnVF6VyH+w8HmyhAAi
cn42dy7vNthRJ4udwocJS/u/OJgqcH0emKnCPtfspb7FX9GIyXomShCegjDsu17D
lwmYKaqJ3kk+B2rTgMnsaPwf24VajPgmMiaTVAdoRYhNLhOzMSX0pzA/gHisi5B8
0wT/+Nom0abqeWgll1kZXufsAqiLONCsBzqaBNTiXv24eJ/+FyoXK13iErp4jADD
Z9Tz9pJCYY7nl7fsivARqTp7sFA+uUIm0YP0EH/7GbXYPxJcg12DO8ljADrBqZDQ
m5ok/ckugy7/qdzieS6LWWriYwHzEa19uI58Xw6+esjEdH+aYv88yYl5N/wUlfR8
SxXtF/lUQnHU/iUVErG8uVDQE1O8plOTo/D8s/PzXyc6c6PkR1ubv4Oq6g2cJpl5
25U7Jl/dsyOAN85NMSVJeXndJxUUXAvvx2eRuYlQEjAqZfiN2UignnXRE45sPtFs
O/kevcsWVOEHBmtr+u1NcdcgcvdDKsT28TX/6G2WjbgvmoAVw5aFU0jmzDHseanw
S4KdFdeVAs1gjgSVK2EPwCo4ysrpVsBcuaRzTgLB2CphPFptgVIkYZLvs/lsp4ru
sSXn8qFe4fGvh/H4u9VLmG2TNYSapnR4BWepi0hV1n7Sb/s9Nm1K0u+T+emm8Yc0
mu5YIS0ynonW80qZPUtQz2s8zcW0T3Le31K8+eInVdp3wj/xKw0PQrCyFKIrfCO4
050GX/Dfv0xSGCarB4KgHKtUe8xYas0VVsQYBWpU6zNmFmTcRqnGgPos+NqmdOTr
uKUDVHNNBU30AWM6eQpbbIhebLQc6MFxBAQe+RTyT0FQIkRXeErSWT7JVwE0Lmb5
DloE60BK03AOICYjYLi00I/DhmvLzQJ+izgMnAJSk3/8zJ49zArkZVgarpeFiRUW
bwO3rA2TIWukAbkASVwL/k8yIbn7PBuASbfmAS+G39E9jlje3OB1N83OIBdPmY22
ytioKSTmxF0Eva/pPJqD0lMNy8mMYzrDPzJQCymS+QcmL9UmBBHt+Ldv9GSJYMBZ
S1+bVhs8/I6QNyiQlhvgku/Swx0VnVwDx4BoypdxT2DTT2zZCG8mjZsl4R7KD+vk
Ezq1OvSWxcVSiO4MUZGU2C8k03Gg+x5Z4scgih70plQtTeBPR1JiW6i2Qh7aH/0E
nmr0fEabcjzXAo8XcjVKjxU87/mj1ufviyy1Imc7pcdZVm7+b/bB4YpdMkT8MgBR
J4SRxa3+8d+UJWPO74fvlCXieUsj4gXwTkJRHXf9/6VZyVbwpsk44cTXsehn9StO
OdZ58PoKMZH9zlKKu1ljy5JGQCH8pizahVJodmvd256cPIALARrLiUjlUxSh2zvd
wmsarf+qHRK9z1iod2bASl7EvPdcIfotf/xCLsZ9NtdPOKbuHdmP7qVlXVXTaFto
9umcGWAaknNVWDIVZPfHGCKFdNhAvEFhDAMwS7b7HAbj6pmCjwhFoupxdNPkmoUr
BO4OKX9qTnKChyLFBgmlu3x2y7GbnVYpmOpJThQuluJm3r+jzLiN/jcE+Xj6f3Py
omZ/hr0WpPpbOWapZO3kfn8VGUl6o6EHGoDrIzlNHWrfROAqYK3CXDJ0JzvF2C4p
hTNadSWt4c55pr4Qrw6ydww6utfS6vUPRCqeWkn92fxXBBBVwV28b3yX/AqVX0Wi
EtoPiv9+ZI/deoGZcCL267qOoSW6k4TUQixe3lIE3Q6Sn7eNpws9qqCRAsk17Gv/
vSEl4x91IxLFwriH3GAJPvjjK7wAHFAsYrVLvjIzIbRCEUx/nosGG7PJSc9IBK8G
nO2W0JWNyHGv9XA3tPqmQXdMG2Ws2qvJlnCfE4YbM82HAeXmkLirg4/zkLNJREZ5
1Me/dQ+MxpFKFikZiRUYIH5qM0rfEXGqj+weXuDdBNo27YE+BDxDPgo7DO6E4Eqh
Txw5MaKutjvdbQmCGOeeNra8GaxSeDy9YYChOD+IEPWbzgxXRYBsIbPffaPfLiqL
kEzEg2vYfWxq7xWfV22WfCPC6Cuj2TxjpXJgqiq/QrVvVzpzI7E2r8sqW3jsPhqt
R5z5Re/bu1jVcNc8kDbSghLjp5OAD99/Ezwltw+aQFKc3TG3pfTGfmndTcAAw7Ew
wQN4pfEWulkbAyzFaao9+U5vu/+B10tIL/COKRmsXoBxyqnVWP1H+caTiDV95YI1
V6xbRbmCYNcriXVwcxYR3ge8/LWk8AX1Fp2ZC0sbBav1NRgQFAasAIcz7LNtmean
1i5PO3PnV6S7Kn46QZfkFdgkSBHga1bWgQQv2MqT9OhLbJWxbiw9u2DppHH9/wQJ
gYR7pGZ7i6nwdHwQu68/Ek2Xwe190E6qsp7PD4CeaU+egL0dvVS12pmXIOC+1M/L
iAeuNhZi7zUFbckK/6gcMmf7bKbW1jilFem6CPhDfixToL428ovavzJ5tQKNaax8
kAl66fMXLQjXKZOfr7dreGNAHPtq9piNKPv7axm8dNbGzQ4ZXv49x3jGkod/PwNA
lVq+iMa73y8FeSnJdmR1rWa+7shHcxF96WzfouQRaxRBnPkAzH2T5zTQnzJjFCEH
gftkyE6LcMLlTIw+2r49y6o8uyCezKsfhH1NZl8Pk7W38mkUxjUiBu1VmROuHv2W
o0iPsH7GxkbS+nmE4V+EMNWa6V/py+l3MVVXSBsvEyWa0slhGuhlhY0ZTaFeKzsi
fQczCyQxDteLX7O67T54zrPEGQuelPu/k29HJIhe80kZRUzaUKOgGcTMvnClfzxJ
4HRyOSIW1eiCcGtovduCcWnMEeBHxqCV2SB8ZNgZPLfyN5nAmZy7UCI2Vbb0quj7
mLDBJmmpbrBFLnck3tGDhZKFt9GoAils4Hqeib0SRgsQb8V1K9E47kVWRweU4lTF
xnIxe3uBBcyJ/LPXsMjXfYcFoPNAOmkgkyLRHXjCsId3M3itoq/Dbr5i3eskOsR+
sZJ8wsVN9mxdXKzj1iY8paw+UmEbzwaofebjTK/Y4CYPud+rTr1OEmUci92tQvZD
zT6X0XbUs8oHnooo1mJy2eEKr6qqmCE+X08x5l2HfF/dqUdyVEAbk7KKa8KT9qlc
zFcN6SFDNOMYO92bdj4T5c2NzM4Of7Yi09fe36HUahMC5wAjqiMka+D46KnX1Mvl
ptlshKLZoADbSC1aUoV9u1hJ/NU82Q07MQ/GoTaqQGT/9OGmIdx/A5YzFsXuY+zC
l30rX4DCfgVW5duWTq571C2fm9ByQ7V9skGXgOdI+6BKcksBoxnxgfhHSL9CiO5P
xP/LImZVZIlg0gTfHMaoarmEM5hNEl+hQ5PUtIJ5oBFTrbcd9qea6g1ecNmcQRBU
xbN9NkmKMmH0p+Z2HoDq/igfTkQ/6qFExrm4FecU2mhGUQ+E0XycwhoOdzFoF5lq
MvwE9LMpEjmETza11G2BwG4kwu+2idVzUYmOZRBmtsuPZ5KmFaOcJNf27ZhJ7USq
w6dmlIMYKLqAkiwMRW328anDCjtPqxM0PiJtJukaZ6jM3lpvYtX8CmsVu47wTbqU
oGTGH5Ebk9SPcPfZL4u5nYOpzc0nB4RTsU6oNxezH2bjwQaWjNLAwi9MzWiZytUN
MNy3j4ZXdRtP+glzO51PsWPfN1OeSswksBRZi3oDs+r6W7G+ubeyO+cs4T7It76b
G9oWtUB9lzokPCr7tgBBqKWkyRLC2RhFBPsleLikHWf7gO8gkE8ZdxHkReXeDi5u
z7R5Zr3+PWsGS8oyWRWrKfHSlCHDw/Mf/J0KzO8W2jXuqa9hXU6FHSYp1MgzYCbS
G9SgAnS63e4IWvi7BjKzhrRzfiI0wgMvae0vzdcBTVZghP5KOQwc268BwRQXkRkD
ADtQ7LfMWHKa7E8kzO7PXCxLE3ZR48scjz2pqFBu4jVtGUbgcIPhFVDedFMwPej4
cLxjyifUKSzhFnP6qN44iqDHAmfPG+k7mwcFw6u7uVtMUDSR2/wTVAeOP8I8ir81
fV0Zk+jkCgeMok0yxPyK2zDxcvdN+IcGpmaIZ35Is+NOwKLSKTGsDgpoOMpjvK0v
AAbAcLt/ML7vpkYVrCt2BJcHBWVz24btd5lnwI3343AU4yPg3dfbCqBd3qcCpF9a
RCqdMjq2ZWKBk+zLg8wmc0sGQq2uw3ysNSjvnbP4exCO7opE5bFbifUACmI71EJU
aphx4kdC3LSPWOw5q1M+TYIF64ELfugj9R784BCyDZuS93olK1tP4G1ohXuutXAA
UUll7pf7h4v8D75lNTGLNKBm5B5TGyyj8/HQxlMAOkAHGJdJPNtDrvQ4fq5wUmet
IaEtRQE9JbOyJPX+aBTJy2YsFt7hp1z8y1sFBWVIc49UJJCzvydHIhUN9iS1sc8q
hOpBT+iubsaeEOk2+9h9SskcWfMItGRAptuqoeHY6C0GbFPAwwuOMuBCRcmrjJ3n
NUIR49KSsHf9DXU/h8J2M3tRvnSMimg3k0LSmc1KPoDEnMssGKUDPJjSP+vLdRoK
X4sgE3wB+bhyfIoqFAyZ0vGRSrTZi1aokidIW/um6L0+Ucy57LK9UuO/4scb5/hz
FF2WY1jEmGnxwiyaqiR9AYUkqaG81xaTTQtfbqUr60fZYWJaloyo7t/Aa4CqnIjL
iQssnNeMPbmmMFvQ3dBbixHFfkJTXgS8n6UN1sa8BdXoRukDj2gxx/5YO1vCMiVl
ASZYtILIopBZQ+qC+gXTCahNAONyRk6Z7vtA8sfkKEDAROOv1TkrqSsmlDAjmcFe
MQAIBfuoiKB+VL2cMgBjxquG5vZLVfIxfAyTw1X3DivjyjsG4WWsUgl9RUbr1KKw
UwSDOIAaFMdMWJueqeQlHgl8VD0aZkmrC3i5wLW+95Mga5OsioHvqynG3ydx+0ub
WXzLD+AQoA/srB124wFc0UPRCEv3QOYvk0Va/we+Y2X/ij3K/6WsthjAz6nljRMi
UU6ylIHfI1tgAAfDOZeGrO0RRF9fzCsMHcTymsnrNIrV/5knyOT58EFrbwUrtwEc
SLog/JIxiLktkiTbqFElvhfEe3/dyGrk5YsjoAlciQUOf1mHR9ftmGCLUADSL3CF
M9f302W/xTYw7oR3qDQRg+d64ch+J0hI6OZrlV1mBIpZuFDWlBpZ8n5GGDjWYiEM
72fxapRfZc77VAe9cBYc3vEIQ4mEdyB08t758HgLtxrWdWqQgZxSbzs97+m8F7wY
a3Jr/pH2YEq5clS14QHzn4t9wISQOfmjPAgNC9MRgP8l41uwFnvQPxToxRFUv+ic
M45/A2a5iQPdmEYuXBlFuTkUCYOTTKapvijqC4QxnP9dEzkOYYGwlb23q9etUaTP
JtoFWQw47fnnB2tbljPGDoXvAKD138x0T/Rb6Yr62psiGZXutnmdz6NVN9YMuVwY
aYl9iKSwjYrWUeZArDvRjsRPJHyK9cyvqh+jIGqGg8XctKrhSqse+J3L7T7ZKV5l
DoQzns0J/WVkQbssFgIndFelqTYNeX01DQ++2nQ2PpT6iEbj3RJ7GdLug2ltCTe3
KsaAf1wFJ1UE0YBA1fPKoG1j3oHqDg9X8t+CjlI0UWNVpaGKC0mmQgQQE149KB+H
11WzO+B3DITZidbQQLpZ587HMH3gkSUEecan6zS2bDtoVUdkJUiwBy2s+iSVl8Xb
lulxJzO31Z9yT7XwXpSI4lnUr+TWn5dRkBWZ+kUXs91JapsjZWQUbCcPDCHS00oV
cOZg7pSytV83VDr1iAu03VRGa4kKaJmqiEiPPkh+3Vj7/pq2A6JvLKmuqpFeoLv+
3I+9Z+OFZORo4InD5jup57dzQuUNERwzzxoNQlWzzl7/HUzxm5BXe6Yg234SwOb8
R20dBNeyEENVnNcTmmn+6fDdKmT8220iAyAaEnGgV7CbNBZpqYwpjrJ+nT3aBzVh
MZUPkjPimz5XHXRfgjSVW8PGpwRuyOLbixdXqHGlmA3jwYe62IDhMasyS1M5HOM7
fbaJHLlKdK6Kdbex/AvOvxTpdXRwopRaL3t51vdxr4quE1IYbiRYJk1R+mThrCOV
9M2DFNCUTcA8/ydVNrS9it1EID5dLjYt7zMaGUqgoMww0/379swQF5BggEIyUOI7
7aRbjZqbLmJl+6vhKacGl6/LKV1iWhlGzIvImoQecdPdtA8C54jWnFRAi8Z1LKYP
1NN3sxPeCz9kfA3ij0cCOCLz2lgmxUH9GIdVZe8VStIU+3rX3b0PAmFtZiKS0AMr
pMsE+EeXLYlz8vAtS2ABfIu3qVGbmkBszwE7Y+s9kjhKnyJxY8aY6EdJ353p4fwN
L42WEIjkJ0mWwooP3hAUrNaKLkQTxNy1Wbhyutitysye97YcQGYNYaCTUGt9joSr
g+IvWvA2YPj7MtRf9uSjGnweP+vOj5Js74D2h4wcGj0bPiZhzi3eZLx3UwqG97Wi
KOQV23wxrMVKpoa+nj3WlRX+VdJAKCQ/4oYCsDwnykV/3Moqvhr0Ckprx6WWAIsg
SqZBHIEvfcxt/aDfXJXi9b4k9DsMGxHzlyVhKtpnYviqbM6f1YAXSBBxrCmFh+nZ
Hb42XGJol/btSHbpNR65KYrMiHGgL0AxrO+DyeKww6H0tgwwXsq7CvwM0Mrysnqx
9efPcyhKtiB76L4HgdZASzhbeEsQOIrUCT/LhZQ8NqyR3amqngOek5v+0fnJDdh3
76sYmc7VQKQNiBRK1ei1ptult+RZsGEjO2Vm8KHZpe3hJc7NV8WLR0dd02NJsFLA
/zZWwZUm+bPGycImjjGBWMi8yeKiEqB6k5v6hWIaqzLZr0zQZUYSk2NaqTjW6Tiy
9yP8n1Fgx4CHNSJfhZ/HwoDh3yJUetDeb0QYNF0IPkrNnKEm20+Q+pMcnYj8ofzA
Bnry1mEMgsbyp2/Bt+W/Tokd0OgV91cBIBn8t4ScC+PAgsapo3fif4qdObRXQf6L
ME604EyJiQyf134ERytaYNWFSqAcvyr05+msY4lJAJrs+IfExCWzJu0dmrtV272k
8rufQHZXHz6Juu68d5gSktqD7mGb7PJTDELMJ915J6wIDW+/BO+rrNBFszj18kfZ
8p3VWhWd/NtzZ2/kqbPMWkFjym5R85M/cc2uM92Wxl0qmulnMyBXn6tReg67PYkp
fEln41HYOANQHcx5Y9fYcWvPEYV62RTpOjaEvEFv3yg1J9BLa9kQ4dWZ2u6W4flA
8hnyQhQe5HXCzEfZd8jbjoDmavJRLzXm3BsuvXvRVDjei4it5ljTZcUV2l/qkGr3
77KJX4ivNKFqrhhXeBWtBbPYEmUnZdMYPOPrOmtMkJV8j5SCN8UIoasX0GQPxA4o
J9vT7uJ7SwN9f23lHuKnDkQwak23v4GCCEzve9kvudYyP8hmemronNeV3htJVymy
OzCMgg37RSiUvK8Lkgt0xBRXnX5Kt5HayI4SswFa8HrkvuK/F5dfGCAYjlLeoGm9
tJ/vZxop0tz3tUiXt34gy8iPc5e5d0wovZOLl2ZTHQi4V6C63Tego9BPChpL8Oif
jhb4Y6Wrv6bfpnvG16OHFmUvCKSlNAKMRlVuKCK626bTn8MgaoW89ajmh2z1iLyh
k5zcZXP4FzSp1sVUlKI5/qqUEc3+OY3K0lpBOH9molTcJ3qqXPHNJxpj+lVz4a7/
GFuEyD1I/jt6ZUbiP9hQGlKjgSCZaZIwiTk1ve9GfRtIVdNZ5NoBkgT4hRrEvuI3
t6gLL4t4alOkZfZPuS//pwI5Bhdp/rWwXRdET4nCrQUxSQgeV/joUO8CQAygxzj9
SSUlDlJNTVNWqlp1rENZQA3IXlXZE/XIVA+Jw90Iz7nUfDUWAIff181dblri4vqV
U+alMP5iXC+w2DAwYjun115MoDHIfYrxxvw2V+6bN57HD7+r6gpNrMxU3SRX8wkt
3+rE9huWq6ElX67/WLIeQwnEGiPBJnWpWWjHU0/u+W0pR+nxQvQeLTSsFhPatyTo
LDN2LxZ89vydtRtjZPQMCGP/Wps5k1ADCAFEDPmX+8SgomwQAxpiKTDqgcu5uaLJ
h1ZjxFWKWBYezs1Mio8ua3Mz1KvqbuhBcWXrVXL/IwCfSe6E/k/BG02lVBym6Gq8
1ox0ZjPooZykvuyXwUzqM8NqV8KJTLzROsxej2k76bea2EsIvOk+d4ycVu4CC3XX
n2wmsmvJRsbISGHBGyAN8jhIeM+SmjHghEcdZEDjntvoG6hUSS8TVFk+GUbCLH5A
2ULY7f/L1r4pEKq4ZH2H+4nbAGCqLNNhBqhzkHI42ZZnpIpFp7KKt9e8t0OXZurU
kpOLj00N+K68/XWOuxSFMqrm4XcNlIxk3zoigdL7bz5c3pUjODPpD8+MYOoNe9fC
NrUuEdMloTSmeQN1gbBMUow1mHxqOpcup3hye1XKNIKYwIhks4qXeqPBhyj1bMtd
lDviEkYMue17rSo6EegfGtpxH9w/uWWbfvoWfkirjqxN8DtMTwH4pH6JOceIGjHv
DoGvxqL3ql8xvgH2hXIna0IWLZG6plTpthWzcFLIxzAvJ7sdiNJoDaFbU+X4eWqy
gAaJ8DLoDGJ6cLpIeV//PJzyXTGMXHOV1DMd8F0i6sTzqGRs+j5ltKVlTon7NhGC
svH+v+U8EjEBAUG+NfIVHilqsybOIg6y6GkeTwOjx/KnxtxVx/9qma6fHSFWJIHy
i/c3hIEpvog/8YaSo2Y7l5y8vMzhDADEzgxkSJFwBoxvM8B+lR0pi2AJ/kXSJmy/
F9hPYeIdaGKPwyCTVcFA511mwN0Fy3omdjJ9v1vwVu+GHa0AoVpWfw0JWPe6v07z
tY+TH8I1iS7yvxtjSuTbdBDEFt9c7uNmB2sFTubkGxfllTPkJcteXHwbUcSKS3kG
oPzm6bjx/0rbSVJNBZJtWwpmhYQYg4JQFK41fIt5MkpIovJeY3Px3SvDqB/DXhHb
kr9ZqAlkjmmTCvD8ycTxo30rid41goVM6AhGQLepC//JMpy8Sa3+Yry3+1YF7dCR
bHcIIrrNgUMj52XCivkSCUZS1rtiU+oalnk0dP4Eg2p+/hzKsuRMcR8J0B+Pnpv3
hxKvnaF7jh4G2FQBKdKlZr/wgVueTD0bJ8zMEpKxWtujVP+ob3OK6cUK3ru0UflO
5OqSnngCBfVmPE585tzksb+sFvWPIG7tlzbrNzdZ3JlHOMkFqRMW6nrIX0cqh8y1
1S249c3xGvuG85ZxPuvV7oQDLVqTqOm7+ijeHAj7i35vZC9LZQrGDDuXGG0AVaVS
5qYy6373Heutn7J7if+UErEk3sFD9WdZTr5mnomaRMbUQSzWXHBC8tUlKPkjjjQ6
/WN69DnMhFnX7SqxK4asEDbO1PnjmtalbPhCRZoK6hRc0/GW82LiAiG40LRYUwZW
CQbQGGYJZNnwnoOMoqpVZH69cvy9lu5zjStRxxVcuLpmnDrBwFA8GOV503rdGEc6
8XW1FsgQtUXLEJxkQ2OA5CONCFgNiUodsi7wsRL0eSkLLtBijms8LcCZdewPB2n3
/RmelkLC9v+nNveS9Al2A43D94nBLat00eUSJsEtUjQlFZ7M4Tl/m0Itz/Zw2ffO
wi7uXL1IhbHqJj+R5aO+0l4MrxH3YSevdCc8WWH/VUXE8tj7IH49+ewQzJSNhMlI
8oOMpZnFUQGxbkQPrxpo3yxcKqoGkd+Y3Be39Ge3UpHtDH6lGzEhvVOcixuDhCyQ
WhPTAOu216kPCX7//1MP2m2vn7f+DLVdQe0Vax+TQkPGJ7hS1IO3bbyrWvFwZEwZ
We33r84KIVQ+mMXH5qVIhYKQrdTGC9eCJ7dGme5Cg1ANYd4Quw46oUJg4Hd8VMx0
9BjvXTEbI2UA2w+T/1shgbiB/9bocXm8xed13cQVmhlYaNCJs4fjZ8B1I0MDBfUX
WuyKEwUtOAncCrZ31BFCD0xP/dyeqpfgjaW6lf3mlORoVTkDXkQ7dYZOCdTyw74S
YHDmqgLsPnzevCFn/J8lJKgTJ5wbKz+ihynkYiASIphprBXpCVTLwbWzKC1uzlZj
F6vkTvrZa1zTbpCvDxvGJ5XLEz4ibFon+Ae/y0iKq0GHzARY5weYAogPUdMne2pB
ZGTb9wtOxvNrwnnzPPLE2hOjCl26RAzAkDyN4AgooI4EAxGtSOtNoWHjxdVt6ZwD
7yLOxKkMX1XgwwvBwUJ6q8kFzHg3Ww/sYgQQFk3ILt6Kel1r+irygdXC8kraliB+
qdItcoxViLAEFNNUogT7Zabzha2m+KtXdrUAElJoWVfkqCGIaQmWKERrgFm8X05y
vn7Az82hkoxFH0gkk7CIXabobnbS4DVumQayFUDGbPy3bJC/KcUgW3wfQOjde+NK
FjYOjAOoVq2Fi38SSe/ie9nsiUOks7YZQSDVk4vOgnYDyCRFxTCOXR0s8xlpxgaZ
IaaCxq1ZuNp1TFBgcFfvEBXN3vdhnktd/CNwZtyX96HeDCbqWOMY58FawXZT6tEv
Ikh3Z0oQ8hF1X6n8eq8A1iI0YlOTh5Z4z5DN9FSzo7+ePyz1TnFPetnivOCXlazQ
ApFMluv2PaCg6PmOmm+1D4L7jnRgNVUL8qyUS53yRTwXU55UfFpp99oQkIkprIRv
+PaPkFUmxN3GvaWQSQCwo8WYPs75H+o9wXAwAsTkS9X7ohVZ5jQPyAeJ7zXoqOUF
mEGUGmPYvScDaeoC00aoWqPQRjxWrDSv5JnZLEeTxLD7oWiMYIufegNb/O6jVckd
Ql/RCoQi2qeN/vM+cmRIxs5TPm2DP+jX8xT5DMDRUZYn6EAsCda+Pre5po1RneUC
/kDgOLVWBLV0mr9JPEB4gumkkn/KCBoxfzDKXLRPeFxPauo3ENEk8YTCuepLCU1R
iCfkyMcAoQZ3iFozs7K5KJ11H04QRD79AULJvX60zXBgmCnit7VwIUvWPt7OlWW3
Iyx6wNC1R6C455Y9tzLqJhJP7HjDrZ3snykit8+L6E3pWLNBH5DxwODzgYlKQRnp
D9+OsLzi7WvymrqKJ46I0B1h4jk+L6+FFlvNrSXgniysQGOifJoNyJMpBjL4vJdH
X1Eh3qbBB6Yimn5t5JaCa8RVLDlbAaeeC8OHGlzTbqgbVQfuO7HZdJmN+Agpm3Pc
LYJAvU05Q7tQx+5bpjIN0ZIPqcMJqk3CR1B83+lnStJAV75HN8m/AZesyn6ljOmf
65GXpE0MuOBjCtnYK6FKFOgZT6jklc8rufVljGFPkCMxdsxzeafXMJ+E0pvI292G
Nm+SD4zHNc8UsIxwZkiHTj6LCFcZ8e28nmypVsPi2PDZDVmA9Ww8IqL1tCQWOjLo
otSpy9IhcPrJnTrlSAvA3HkN8Xyq8OI+qu2FpNTYqshRZGFTy7fhUU0YVL1tKKao
okXAp+N5nzVoKr/Gxo88L3ebebwFG4qFTheW6Nn6MdvwRK7clefZ9enAgiXSi+hV
njggh4pvUYmPU3ReyofCo0rQXieaVi81xSLzuG2M6JnG2Zsu57kYYO2VJTPkaxFk
IIjOVHZukIaTA+ciJ7TohacktQD13eOhz3Fw1ad/OIGYQOWcYDXeczORdmBCm2yH
OgxdQOb1EacU22vdhmxcTMZ4PSqYGvAVcInoBoZTf4MgGsFCu/KqPx8B1l4SRVC0
tUgcj4+MWg6xS1EL/cL1pVaW+NOqOCXN/FQrLQcJIZGr+haZixRrlzW753dDHm33
QuJZEqwpDq4Wt129VEgVPpVPnRhMKMemQMuoFfuoQLo9k6evCHbgiRBNiQsBS+/x
GQ3UFXUz9alYBIuNMK2lH5/LvVXIzueTc3QHq3smzwFcLqVpukvwAAtibL8cm7ed
nxDq89WghbRUr8Adll3HNEnmaXiAwM/9k1DHG+DQAOnXiogOYP4YjAkhROdlVLBT
Akzmi2YpdJyC8wDff59iacbEsBHWyHOpX1qa5pZXDZL8XiwSJfNoQGmumxA/87R3
ueU4Ri110sRX70RTJkIT38ZY512uMJulkw3SaDmpXYNbwcJNowu1wM/dykdnYNqP
bnFtILekQM3k5pqEyJbWBT1QvHYI2Ugr9zH80lIBBQpY5Spm2WapSHb0zuP2IXDh
Gq/+4Z10HPcKr+ATHC5L4Q5mUvvrMU0P4V8XvGu2pISgSi4YyrLc9Ykn9AU7SPjC
kjKYrKgZs/HHoTJZsHAIG5hwEE9g2MIM2coMBahz7hMOSIR1zPy7WRBNDO3H1bA6
NzTOwS1q+/PvJUKxAhA9LX7B5gQT7oNA91YPnK8A+4WcNPcSedJaG19thHj4foR3
pI2VntBwiItIkZAMQV1EbJhV7aJXvhpirxE8eihidUfubvO7ZQbALrfee3INeUTM
CyghOfaaH6l77m6dLFp+3ziMVvZrKa0r2Yr5UJDd3+OWxaXv1V2Bf9Mei10Pt15u
DPyYX+QqWZZuzLZDUtb7KZVSgdr2Ems9ZfXhxkBoGKi6Hb/UZjOmtkuZ3Y/nTgvx
XeLnbg+Bp/PWanbJOEkm6hKop93xB+RxiBFlKa749qPRSwCZEbHlp8vlKfwkw27N
0of7/0wZWQaFsfoGwwPfIPOkpKlE5X7yjtmJMAAC1m5c7S29QLtHu6XVnMUcVp5L
wPCYpUIRt85kKgJtl/PyS8xc0+alHUqyYtDEsSX7+TCAAjjHRjgZSz3tclPZ5Fnh
UvW1Rr6O19F3yM4Qj9gp2XGX4kjPb7NIeOk0KzqGYTvjK1BnI2GmvQu8JEP0/tEb
vvSatGm8Iu6tP/m8V8wkky9y41mJ4ZJHhgg3gHTG2cum+yPzUvWOOqYgu/VLMBBG
MZfQ3ERvSeZuf7wq1JiRDpAz+kaf9A3cx3BcKISxkMH9a6Hm9VRdJigCWMdR2730
lf46doNiUt+bFHt7iH6h+NwNd+2EwEUjcnTxCr4taDHBlFvK3q9fkt7R3LxGdzdc
rKBV87ST8crC6QIkVULbL/zwCDLcZaQ6rKCbdzGZpAxVcFdCCggD6f7j+nfQCq6o
ToPx7+WV3NLkql85kjzR8agYdTrsTQXUfqtA27XzCfD9mUgGB0f6mrAgCipDUlhW
9qOOQTJQm39FdhL/4HLUrqpvl5OH7Yu/OLdVfp9p+6Bf+JCdoO9Dm/MyUaW/DTe2
FUU2D+MzCocmV8yyjz7JRJDnEWsFwCB19FV0g2I7ndwr330eOYqU9772myiPGr16
qi6x/K4hJMNQXwrSL36cRcCAwIJ65fAc4iWVj+STPORZjtuAm7Mdr7wstUoS9y4u
EIQ9x+GLrwkdyPulPknPZadxUkh//GR5uYKD/YTFawT/ocueAihfxJG098KsIlwP
QsANA4GttB7lVpZCwQWmyqg4z4NCSZ0MbFTQ2EzuZUhf5T+puC7uUyH4pwQRrwW8
G0qblEdV3zpWQy4vMQnJNHq84UX1moawLYBDxs7m9KB30qRWverslVlNgOXTuJBJ
RiUu9N3iF+6FipL2qzXlC2lEQ5Dq2wvwdE1Zkgqk8/AqtT7s2BmFXXFVI3d8twJc
SttEUpnMopeK6P+1EfNJE8A2ka4tpaw91VFEl6Lp5MAJLThYpK1jnSQw6AwYN8Q5
FW9c0Of5aMIsaqynlmD13uNr3tLVpzck4ZaSJc5a7JQOtRJNw89LuP0fipaR1gyx
0vFisT+8BcybhVnR1PjP56L03t/h4U3PdkRXbv+otLT4ZF9PNrMSE1AwdU7KH1Il
NNJyLBXtOnTabZuiIlnUCiPKh90x21v1s1EGVp7rGANiYgr+qGiM/xSnW3F0SD8T
8kptH6kvGI3/+ToFDnlcH2ZBBB46Q1lbBOXq2bXROREX/fb2e8querXqnYwSc3H6
z8fY2qR5UKnfXe00zgzfeJ/fm2oJlz9KBPtrSGx9T6LlFuU7PzSZc0gMzAmS8ij6
NdlnJXPsSZ1owWcyk67k+UB2jO/y7TTnMBmi+24tKCTchF7U6B8KuY4cP/weg0GV
U5bIOtUk221WnfUFL/rVE1UgCTKWgat9GjYNtss1OTln2UNX+ugKIEuC/+NR1XDz
u9/1fYmdAnRRUPdEecoknaxkndOI9r3+Uwts/hdtRJWb37iJ9+XVcjdi2BQbc99v
nyyh4aN++eXg+FkNo9865IYOozZ/ajsACQ/5fXiUdhfvKz3usdzAJdAa8Bf+m7Mp
4drnKl8qUBtAKyxYCbr/1HuFmQacLwLNkeb/AeXk7Tya+CaAqaUnefFkTd+QO/8q
jwb2/BS0M6Archq9LPFt8h+uIJ6Xk+JJy91OsOGy/FGLvLKOnKPwk5KGsUrgQaHI
S0tfmJOwBbKd2yp6/L3KIGOm4rRiOOfGZqr/yGEW/Ywly9UNhlew+AfWaxXsZNyY
XmeXOjvuz9IJXmBkc/HeCDAGUkor8S23NkleJziQeIYpmglPOnb2HfjmB+dGPayO
AWVGjHiQcwd2ZVO5GJHYFva9qlcgCMSYrKnakEU9pW24Puss0JpEXJJ1W5qJIMnu
PDsBZ09UxHTLUficcRiOfG98LpuW8CcwVbk5ifJNkDDllg9VQr8+uG8f2SX1in+/
kn95+qyCZR22OW6QF7pRlbYnARSCm81eDPe9mGKS52qy8bJT3Cnbdpy4noFNAd6C
2329yoAz6BGDIiycN31BWTir5KCN5V7aYO3PkdndyKRx7mb0LB6+BS8hSsuDRLKi
MJeWatpkn9RerS/9EMWfl1h7Acy8UjF80dZbhrSZ8d9/aMKU4lHkSNcI8BBB5CUo
I5XId3wLjKdVBuj2un+WR1P0azKqq8w5PmTIOLB0R3/KIN2li87rlSbeX9/WmRiD
dUNfvFJmal3ds5F9PIYOn0aw6Xlk2EaWLRcXsZDP2rTIj60N3434HF4Em022nnpj
Guh+D2iDgfF7rsmaHixf8F5f2MiPdF66OHYUhVeL7RZfpAH4Idg9LrOMnEVqJ+zu
iy9rCcwtVhU54TJToHT5rRZ6k6aROnLVtfX9/EtTT/rSf6FxDhb0lUJtIkyvCohB
vLW73M50v8sZ2Lj72pd2u7eHs1YhYBxQhSkraDiOtDYjAOt+iQLpo+2OtAv3ANsA
Q22PgfTh72Vimq11HiNDrSn99zPVOXyielxCzsD/qI3EJ4G+lVHyFoBNPBsNPN7G
D6xvTsPdSAT5t74M4j5CjWFuRd2XYr+WDkmhy+HV4dKjAM2MfbAYeEEwx4OFbRuD
6JZVdFgzcydr/W7OTNF0Yle2ZTcEzvTaSiLfur8qCGpEKzjej16ynEAk0DA923nQ
/Jx5HZ7WywGxmIz9dRT4cTGKcf37l51Dbs0A3bnc/MgJPFuzjUguKujPv6ffqTYc
8teN+DGcAmZK51U04PTrZGgBDD6lTxrXfIznsQPaWfIGfa6I5lMThdVAEnC1aQFw
9Gd6fnSK85L+5tYZroV4PPYkY7eaznbRVCdFhZFHZ0J4XIByokzjhfaeyU0DmTNP
m/1nd/YsQM/XM88aMkBcOzuVA0HpbrYoAAbXa3QQ+i7eOpi01A1hM+BG22gghAiR
s87SucSz7mu496O4iYqGoWFUQ3s4w/eZaS5rV0OnlRBZwiKCTSEcxcP7O15Tv6HF
Spl5BejKLA0VvtDpS108QjTI9Oe6xNUlKgU1HehlJ46lzvrwB68IVZgTUxTTgy9F
PWTvXJNJgvZIBvzve/lN2latkMPt7nrBlkEwRugdgbDaI8/BRPjqPY1h34PkTqZr
sgZ29mRIL/0CwgIWjGjImTyUTRfSAvVXwBIHDHJCr4ftSv/VLnOWE4efih6kZzPY
lBpTbBPPvDMAiMRR9nvYsDwxkYwlH90LUcCBnHJFMVWN0Yz/sc9HP+gsg4gENzNh
cAFIEjeTBK0zNVGduy+AbNHeDhgqfw5u6CHiGxClpcNrVnnBAZ7TITEkswpjKwJm
kokmtohFLxoWffbSj2zeZfnKp768aY+/uXxt8SRgyIyJOeVvkzHacWq6QYUQabno
x0Ys6vw9l6SMN+LRNcCGB3PP4eItCid+b3Q+c396tkR1s93Z95bvQxJ6f9Z1UupK
PSjGeoZWXH/rQLXP+rsuVP9b3HwALomybsMAEbJo7m1uvyFoj96JcBDZC2cWEae2
+fahdFTVqW7LYwZCpOErWT/aFar1bnvh439HbzHz3SGfTGpVHWfvJjnX/cWUFJcI
Iq72SMhqSjqOKHb0FBuF3YcvsjmR44o8ij7hAErqGZ+XSliF0MGWStp9WQhBy53j
H2BCbvFSKTfG9JcyELYdljY9mlnpu9ILJCKnkPm2FakzdIpRkyUQvp6rYQH3xXTI
OdsxmA42kAAvA9H4XFBs/YGYx+WfOw+v6DqlFjZDAvsQbcOwiu0sIoAr25PlYIc3
jLqffEqDgyMQ7Uvunml8Z7v2fKCL6ayLlEEnmdtvBScJowehkp4etIlEp2FGSeFD
9R1asaTOqfL91QVBoMqGgHvqHt6gHZG0B+Pu6ELnAgRyyDk9+4XM75om2JkVLtYe
iGDZKlVlWWPi7JJsNXqSe0fw28CfhXe9kGmLpgvqTKtPIHOYfboACaMRI98HE2Q0
W8A2nxTR0kjNigGhICB2xS6huOyjnq98VfQckERuffdQqZk25vU6CDRd8eP7Q4LM
IeNkSFFAhlhTY9Rt2MVj1iZL3OkWPrDY329RZmO7QCqJNxZc+pWujqHKo6LdBTJm
bXY8RcfLPVdAL4Z9eHU6F0w3HnaGIBUCvZ5wTNgVkSzbABbLPaf5Faqm3SGGfnkR
d3GT5GPN4LyPShqF2nI2z3bTc2u4dpizEoJzb6OfDAs2HZlk3eJ3wwn/67nx/ZYr
PLvhx1mHoPUdknbLtVb+Tm1PxklCrbM1mgOVDECUZnjZpx3g5lgRhRNZzTKSzJE8
L42sAqQIi9W6Nzp17C1DCljrcmqPjRFf1PG1G7nVvqGNV53kfg+ZUkgoJCOXtlx8
ykPfzKR77U2VISbb8U0YA/8SP76YQw2s35wuoR3SRiAsI4IdTGofpY0/zHbSKDMG
xdp45LUxUcyDFr67aaNcD7qcHODSCAdrY+G2afRVgKZJEylUxa2/qhG0YdgFpsYv
khM5K8lEAGwAbn9GE8UBDji3/F91BDdZfwSWyVBkPUKpFJX3kfhHrKaQENACzbGE
XPav2+Kvy98p4+KjPcGTNoClPcrcAY1EOt0VRUSCZqfwq69C/BZIHrg7Z6Ev07zz
G1NbDWzZx1ouFi2js++Xg7syFboBWoboroDL9nESIokNMdxAyfS5FyQyWz/hbHHT
Jh9rEjEHwVPxl2frXMf5Lbn094P0ooLQcRdgqxX+EJdhxz6bsBF0P0y/GvluMZYT
9OwP38uuqUAKsXj8gFOiklZ5y5VAFyNPj0t9M/5KsKQGlyzNyCEaXfscYNmoVqwL
WDXof60K4/wlPT2BL3M7ko/WjZQSpDgFn0lZCJs/5E0SID1jbw/fx9XxVephHnb0
u/U/fB+9Skc4NMJWdgRLOVshVyJ4p/UJ9ZKQ7q0mO9q/Q2T5e4TpTLNTkk282uUK
607HAbf7m4uUNvGNoOjWl1C6aUHU7L/1zjE5DTpFSKoL4WkbmKHyznNL2MIB0JKP
Ha11q/Tklm7o5+r5B0g2MGiy4K8qjxnuol8Q5WULucNmChWqKeeSXOOLci4lxAU5
UtCoy+r/gJ0opDz98w3LS7+IoXW9MOjhp4ku4jobViIj4+DqgLEpy7Tl6zS30u0Q
VMW6Js7oyyQyE2oOSKOsizh3UgkBeQisrhYS7dnmeEge1YDm8//0dLjt7kfvmzoX
zBGAtqUwjuPkiwvMWZNP5LP8V1kprh0bNPmEFW+6IXmyxGThkqmxTIy9bHYodMNV
DvkVkLXCg/g0aUfhYpejElugOq5UKqBL7lIGEBy+7OQ/IkEq8vpqUfHEyUrmYcw3
J6fmUXqdoc9A8rxd26L+clkl+/VZPRwTRopuQ/YGxE5PHNtUYQwyT8DqrEpBzlnM
98Epp5BQXgjjP52ZKCjVvpyg2I1R8Ene9SRTa7laozIC3xdooyS2a+KIP2XwlDmC
vHq5rA4yoKL2x27KDQPRMVpUACu41rlAxkaeDgTHggnwKaRSru1FAm+eq+uIl6Ll
n8PYD29gibsLPuTGQMgvw03razSWzocs9vjngT4PBHe8+ONdju7DmvipoTxql8fY
V/7fSQtvaQgccjSt6t4c7BZqzct2+CzuB6lx/74ZPv7Kxwv4+QJW15Fbg+9T/aMJ
IHuvIGNVKGeGMh9ZKD0htN2Nim1/m6bz6jaNbpASL8CU1oZQu2ALfT3zEkUzw5VQ
f7sUZO7sBr+Jl9z3OljkvifZBeZy4yX/yyjXjX/50vYRzwdNKtJSNimMpJ33QtBG
zstyUkUYuijs7bBUptPbo5IayEcI4bt5dkLrP+9a5o2z8NV1exMpLgaPQ5D5Xb5Z
XWqnH+IPQPM3/dFbPq1P4M5L2zhUoKxfqHmm8IYEYlcGwH+4oWnXN4usKnFXflm5
npI+rnr+2oE93fnl6k4HppDh8q8bSwzGn2e1b9/QwTKd6Wxx1EeYpUw09paDucOz
IUR91iLLWfaEQgJuSpExG/0GG3Z42rHtZhDayHmIaNZUnI9/d0ELiL+v9GqfA8jS
8CEQyadWq1k+HDgLmQ8haQHKF77YU7q4514nQsfk70gSF+wuiWRhXSsIgAg5KQHm
3XX3B0Iy5k1XI11i8/21DIp1/sR0B05GIlIu1EyRkM62Ba5KpSnQfeQj/5uxUbeE
3VQPbUlJ/h8xp7Ge1752n8yd1m9MN3nkuYiEtqz3sqPfDhYvsCw/RbjEpmHdzd/b
kpWrif22xebzvjWjs04EGOL+cF4qDMPYUf8z8ha91HJTUAXfxjYMb118QEiXVOvg
Myfg4V6f6clAmTDAG0fI2GMPle+hJ6gbMDhdHE1x2R4wY4zD39h+XnIZNL1QD4kV
qRAhVngZxResi27h/mU2wWRS9ptu0Jhv4tygkMCFACqcl1Pdrdi33g/iZQUCStSm
T74LipULHltwVXOYBgAj3qSvSOb3/QDtu/rf4gl52xuNQHEsMMZymGxIma+sGKO2
5Q/M1XLEkvbkB10Jw3RLVg1GDpuxnydDn/DY/6RYa69pcPJsOPlauzbF1r3Bakne
736MmlPyTJM8pL8AZRMONtf10KRTkHboAa034tY8bo/rBHRmHlS7JS/sHpkBmaGr
soZKBaVMeNhQ6JFLyc69XxvWCfGYXSmWYLvbuFMtu8l1LYUd+bRWjwsEhIDZuxt9
DBI1GNoenLQD+a2AiOnaKP9rL0h9a5EIdDKHK8snUn3kfByAzx5o2JS8uNZGlYhV
YP3hqGUXZdoX+pTHeG74XITXfyiFHdNkPVCV2zFr46rRoOiH9Bz/SxFPWVazCLLM
bxxpRazjQquL4i339+2J9dSxvAtftnK65fNeu+8reJrzEh9uCjwfZsxoZ6ZotUhB
EFTVVxyYz/DLPsn84YVzIh2Ao75qejeMc7VG5+cY53olRiHvCTjJHMDdeF4TS3ce
bsuLwIAbh9il/EER0lizsHGCMoBYlXLrlImIu6SIoicc3U7nU8jC6lV88/Ud+Ajk
H4AOGOzVLPY02z9JzQIiEH7lhAHfFk5x4r4stgRZ+IJg/2mh3kPYo8IBP90HlgzW
EcLsQmQz2mUSf5tCT7cj/6bvTUEuJ02Q08yf5yJCYVqx9Sl9jfo0U8oJM15dOIXe
MVaYE5s49su12T7Opigw5B+DSZJBilZ99e3qxeFNYjiWWZqdnA153kCAJc7hkr7e
GM9H0EWHVRqkFDId8HivpIPdTPlpfwZojYwTBIyiE2Cf10czJ47hAVzDr1rdtUbq
Vkt4dAEetF5ZyUWHSzBvBrDHthHBhrjyBIZEI0OXPCHGUfPggpYnCOLTvRUcItZ/
A363YtUlh/qkG9F4U4OxVvVa2fRF7+bX6Wsd0clqbBvp7ehxfSSchadVVhNTQAkD
zsnjgVuN4hIqTmGwVvgppiuciN3tdnOOjG/JiORHJxus95Ck8qFFPypxYEy6ThbP
Ww/MfZw4pQYa/N7/E92zFuhr+K/O+bIr/aXXplUb4dNaTL1f8haR9cui2dQgXYRJ
rveIzo6l72vuQ/o+HdbNUGld60sHNX8FtnnXpTmfpfluJFKVN2gVB+LDSnPOHjKs
jTDwMelGP/mjJgPsP3pdN9Mpf8uagjQWHlh/NThEt7G5eSMCC7J0l4QeBDe9U21y
eqngwm3MisBUECidx5Ych69ZF1Nzw8rrT16I629VAMPV+S6+ipgDeK2X2Jxl8MpP
sW+usGZwGopT07KK433U3TnAs1UtBA1/SNaQ/yHUBgb3jFooNnAE9GJo0HtI4h7o
DlNkkNx3fs1tDQKzVqKB/DHF6rvw7Mdok7WSVB4qer+9jk8umAO2ARr3NRqzIhFm
eL2pfec2GAkUMF9rFtJxf0+rbY2FQoiEynan/rYggN/4gSMEiWimqSUCJnCXt7Eb
70Atu24ZlmIJtM4zCgfx/SHXc9P4QBbMp+8f3XnKNmlrgnjk5R7jDzEM/uH/qj/9
Mmw2AL/JSnVkbM+yHGOj7N32Q+O+FhKM3JVZO0HVwWZMGXBTFAvZC+wC0MtH5R2B
b7utqzrZeF10PjwcEPGR15g5Ah+zEQsY8OE8+xd/FgjEK8bE/qNR+rVw56yJUbQT
QbRzc3SezAhJEa2IlL+4rCCNR2dhlPzdXj+qsVAn0LVy2Lhxar4dphEFs9OrBotR
IEOYTX9T8WmMGFf58jYPSzbV6TDzvy1Di2XxWe41T61YIHFLJsARw7cHigXZix9X
K3K5D57a3xH46zMZblLAzVGaUynQh3uAGRYvW2RtJlMSW9VMGm7kw3Gz2RQu8Qc8
ZLNPsmGaiZZ2UmxW+dS8zwETqwsU2PGMHOeTg3J4YW3Pm2FVmDuA6Sl0Hs5r38KF
xL5x/O2bUO/YzarkYx1VDN3SNSlVda69lSIVJTJOB9n6BW5mWH1TXx5ASOjOeJlH
5GTqw0knHqk92ZA36nSxc+dUboAD/IuUcZglTKxj0V/tIT2j1mAoF9Wtt64/qhSy
sERhDZdO8PEV7D1aBEToSLyNYfNt9ec89Ho3Gc5TZtgGCpZSYP9R1lucJjyoKPDw
dKBXlUZwafM1+CouKwEd+g436BF5Lya+ijrpcnIBteIPS9OTPGY2PV2AIzGsQyX+
RuR/5pXVehlS80MML98M4W9/7zOz9bCRW2hjo9FzSMDaQWHIy8pEH2smwRfpifh1
Vzx4d27G/wc9lQcX149E6ShoDg14tDyFwfojEuHbZW6fdsvzJYFpRMV4RGU//DnP
0rMN3hCnhtSr9yfbKw4C4fVk8DhrOHrCAKWPdmQp5UeeszMcH1PS5Q5OhyyJvEIl
7CByahjNWTNnoQntb0blNdzOV1mK7GSy7jzSP5r5+FYgsj8Q9Selh4I8cSxHUKZe
kS4Snh/4UtFbmqi4gOrBfORddZKPEeDKDCmlTPSDwzijSI8W4rql1i5aVHJgFn7x
wRrlnxE1ZwE2+Um5bGTfhb7Iyoep9K21RI5kqrRfDlqnrbamQQPreYZ6QTRxjMbu
b5QzB0wDOhFf8cpz0OxJKQ1p4r+E4D7HxSChKp4gn2+8FYLvsLd1OSD8rRpb2P+0
lU4HZ/+jefc3O2YV5ahV/66Urw+vJDBVqJwISExE3jR+E217w47RyyHkcjuN6N+g
0RXBg17BQZ2ssXTJ9VZcYbhwX0Kc7iRFu70NwArwe23dnVLY7Gj2W0A5ahURHfMF
DkKL+/8k6zHZpR9l9M7SWwmdmncDQZuGK7gwr1Ly0YnINz43nvRVTAMqf3K7gQuA
CPRhy36cTAU5zrG5jXAin3WUba2QDhCXQbJlvwONBfgBPfD3Lc0CQ2zTtIev8jir
suyBJnyBAAFi1iFFXGBezGfiKC3L95c0KAGOWZ35pQ6/MpkQg3OghBkpUgQ4qIfm
wba7Yaax2St0tyX8aKRWhuvd3Vu7lYt70oajljgcgdbyXGK4R25EOnwPUTk21jh3
gdVFdKsyhlqNf1nkPYRgQ3FJa8s0xOytWl3aXhm1A56CMUgajIfhvx/AbeuMGcg+
CzBqMpLUXN4d8NGGabd2WiTaiwk15nVCP2BvYoaFN2Fcp50rZ2eDa6McL89Ae08R
xsPJUq5hjtmPUCE+nWJ9Yfiof37ZsLqpJDAx6Cy9o4eyKwYSbZwJ4TwebNnf+Zm9
tKnkDrEdcEneoCBfvlAWFsc5TwyKLQX27+RKIYQQn7cM2MM/Dglr7dtaVe+KkB5q
c8u1S3Vq1v2DnlO99ouwWtZzZhySGv8VGbdNUCiQdqF3psuNyVo6rqYh4VgBk3Ul
lfADCGsb/V1Z5YufVuDoZXRNsMt/NkhLbRp6/KH6u1lrz4bGibBxUuoGRUPU9Nbb
DIHY0MGdkcgrjtlVcu1POoK6nWGXmUcb5wepwvboY8zLUUO4GR1MBUFIf0wgAOqQ
oeJp3FBmk9bb9VGKttLTWAWlChp2kUPqKbcucqAZV5c69d4x5KJJO0IHvMI63tg5
5p0o6XUOfJjcJ/LEOqo67Jt8woQrUOi1tRXRgSmEjrmYZck3yJMGAif+SahIiC6N
ALstsG0Lt0+7HuhJFPaZonc22GQeSvEmtkLpGSUexJjcMz2N5UzlehNJFLBRSaiT
5CLaWUBILhnPMu8zUewMODCm0KKEWwqFJNna17MvvgpVsMHq5ncFE9N6ajgOoqMN
bNTxc5Zj87uDtJvWT9lMvqSGYB+XdFlt/4tmPjJNLlnGxmwtQBfRz9yUZd+GzEQw
uO3u176CkmjlCO9ZAi6yp9frrLIKLYStm+QFyqbl9TiXCi77CWPtaZMKnl9A26UL
2nqPQkpSUBIrKdfJPV53Yt4ycI5Y1t83ZYPCmWKfc+EOZ4/jGhwYtDRjFresxHBu
EKWSs/qTsTiGWVVdPXj9mSDToGpYj+0kH8H+PlwEX/Gm1engD71Gdj7AWQ9pjrXa
7qoAUEGz1xy20xG640va7z0Ah0PkvwIeTlYBRbxudBDX2ISdk/V2GaH6wdO4cs/P
DvTgXlThc4wOwqUI3nfgju1JPrUWVcKCb7tS4FXra2xHLx3t3bQIEpLfDVyNZCEz
uCUClZ2GzcEkgzwemuqXnU1ayT9Ie6Fuz7tbxJkDuzHRvcStjC2kq6rmCDgwSFBd
55Yjouq7AoqIV4dsm2LsBL3z17Jxw0hDRgSSv1iv6Dfjx5GpXZWb/yM7lRSx3XlB
/pmhVdDuzAfRswWKezFfsv2ZptFPZUbsoiyZOkPhnKXAUk5BSb/8+hNby9HHjcu5
Maafolp5IEYtgcbGW+Dq9OMmV5283vr3/hz5vm3MmuuELhLz/XpLUSD6Ui3MoOrM
b5L8tIU2gJ4yV8g8iwBGBlFMzMvkc5BA1oQIoK1LWd8yHSuJNPmXidEWqpbONSfP
snyzS02ICI6tLZzZ2HOTol8PZ8USo7OG+BNabAV9ZW7DaiZWKM3w+JMebV+jqFiJ
PCbAleIzcNX8lUlSlNyzrgbAjQgS8kZ+6BLoMiFZJTlpjdll6DIao6P8RJZQSlKr
djjL7XKhBmlUxLbjZl7vqOxQt8Wh/3OLJYHZgkdeloqRGqHizT51KhZw3ixbfafX
ABFYXKTAj0bxmvgJmnkfbzR86s44XjtelDMF83O1IFvhoIx9bdEwUA9Jo3bF4vac
e2CkgutMCbY1FqAAFSqDSZ04VegzcSISiKMBhaospE1+lH0b8XTPwcSElfDX/+Ho
D/nF3PtVFQPqAerhSU5ErJy1rhIV4T6seEBER4aTr6gKae8qc+Hqk6Rdl8GwMbbf
7kkPgxCEfA6NrXhBHPpvV+7m/3vyDe4RajhgaIIMKcDbeYPf5XGx66TeAhvtqDRK
3wHRkVWxi+n8VEkoRTF5KCMn3q722Trm0bUuSk6VdSTRu05FfK2+rEZjP5+DzV9E
YFb2Nn0XTpddZRBXcMtILw4tclF/mPUpmtdrXGsCLU5JI/BfYKfg7NKlH5Dca1H8
kgJ5MSDFvB4G4YHKVY6IdhMk8U6cP7sHt/HRbOKdZ6Yg2DeXrCTmLs5Mx/I1NQOw
TwJxO1To+VknQC4BVIl+1LfR9QItJSuLqzqKKmoeFB/6CjWaqp7pCSdlkNWUIexF
Kb67hEH2EzOuElfMWK/IArkNrnZaLGGDA9alLFSq0STrgMkaIGRFuT4bRcKZCmso
6s/yHiNxN2oMvVF/rYcSbyzd7h+8ZRtqp7ZCbupkt29LW5KiWrIWBqv2lhEebGqs
7WlcynwMtVICy2URoIPZ+U4USM/cAG+WMhbOATUIzV3XtHKk9wOfGKN2sIt5ogCv
lFq5O4zzaMwJ8PLbb8NvquWZibd2ihVVrm96bXAaHiGYMUl4uUlQBKOFTllka54h
1rKhb/0Na9FzUk4BJ+EehYcsABaTSakBi5Vo2uI+XvXuaWTcWAHCko0DV6TlYfNP
lWZIMSvBz4to9tYb+i6Wo9qI+EulUsphJclMupRJD6CqGb2GwS11amArBPEsNSxW
GPMbFy/RVp+ka0Wx4pGg71mQKXcNf9WUHH1KJsK2uPRW1o2lH+v3b+SNlW+mV/vM
TZV9dSti6vje6CX4vApBSS6TsO4iT8Tc35O7UfPcLPMmCvMH5KBxU4OlybNmGJrc
jY6Vf2C4ST2dMDVbvOTFbfB+8ab4HNsvVHGcs8/1G0jFyIL/g23FMo3mLxBj9Hr1
Gb8lH2Ci+w46MbP+gKMIlme8WlNMm+L/jy7hImyIeDpbMMs6W+lA9Iej29GnniK9
l+OIYeW23Racaq8CFz/rk3jvzaF/r+Hliu0/z3KYpN/eUrNN1cwsf0XVYQBzA9C0
epsXkAX8A0ywkI+u0D3WyW1RzFRUvHZONoK8tMmL/mMcDjw+VW/Z9vsTAdN8sP+0
dETLTFE3HNZoht6GItDZ/aLrrMbpNn3rZ43tUvW7dUziMdvDp6ntud/LfMqpVmez
ykE19QSDNwocsiGkoEv7lk42xHuxMiIBI887aKkrBmeUkQ4wsm8fk/zjyawCVkuM
mBh57RH8M7dCOWbZzWcD5ydew9eNZ4WqUOIL3eUB+yIa6QCWFHkBN5NsPkQxl4WY
rm6U6COzlvdxuhlgrZDSC9B14B8cf8/gaNJFDRKdy9DoFnr1Ua72BrpcqdBln2Vm
cuC3V4HslJUrK7s/q6gxfq38e/WwGJPFEzVh2MVc8QEh4QPthj5X4VhX1gA79DOt
S2x5yoCkPj6LrHWT/8Hdt1bgfID5yS+89gKWflfjsc2Ujg8r8VQuu4HaWdmPjTtl
r2AXe4I3sBxg3uVIifXmUbtsOwlonct5kTR3ZYYg2GGsgy27u2OBqhPbx56daLYq
O+xiwCM+Z8PD+zYQeYLizg1k8DCLy8EAaR+QpCMaZHcnxsDUVS/GyFyreFWyETBS
E5CFjnJjyVlnL9jKchFzfSwopGOw3du0APJ6hovS1Df8zfWtCtg8Ta042+nSVU5J
hQcUjwHrkTDCD9sBzu7LnL8RtshVMf9uCfl3xaXJw0smEBKEkwJXR8AR4WF7zjsa
2/qHFNtncb/ps07FSIgwP7nZN4ihJ1e7TljdvOJ4G/zjH5Gbzs6R1k3PIsrDF5tX
mpwj4VJTIvb4ClLF0XLsrOplOPSoBSQmdQuUYy8ytZAzy0ktCxkzH0c9MBz/1nhU
Ciqb9kVSsCktyslfFWEZcYxE8Ak3hpTIDurc2nxUxyUs+xXxD3CUi3wrj64f5Hbl
UVWbLAA585iDT4DlnZRlZSQqRfOMFNO1FgVvqPLzCQJxdMf6arpzUOE2O3zvCqC7
4HJp6Bj624j32Ue0P1xrTRQ0HiJmTo8heynRaHXrkN2W6L3mrSJq0bDGekH9UXb1
nm5diCOSaOnW58pStoUDrENYvOcv3eOq5dXMtFAtVwy2i5U11WAYpsMPP/pvNPkg
HhfXGfE631bKE7eYi5PHjZ0id/ezvIe9GHEgmegPDFaKFGbXqW9CYjsc+yRclmgw
NPWOJRB6nRbqFrcBhpUKj4ZuFQwwgPQUvtlKQDvfq0lNGr6/H1rkrBZOQKxAuaDE
2TX5vWYB+mCYtyj2p6BcjQKB47DGkDA+uRofadOW1DJOXZAGs19fb7m5lywjYJVA
HKZbx3xncjFi4mPRrNuKRywQq22fD0wMGdKodcRnEDV2j5Sfw0fyXBtOoJSe8HkE
dCpt5rJ2mo+S+NBSaIUfd18rj1YDhdZUzAgOUnGCEgpftCQLPxasAGiC8w7NtU4R
MtYqWvMBzAYIP1wK4ggniCLw+fVUMkTZRYtITlZaag349IgX+vk5fnG1kvcGwfUO
u9FiT9PlYvYhgQv3Nq3msWhwTEmOoAFBHgibU3g8k1D5YY0X+Mo7bXwr3QgomDNq
6wdQ7rbj2C3aDikk1NixbqgAp0BpQWpEnwnuM00eSv5MnqeQkIlwEAXiOkwHVNLX
cmH+I6V3xpyAHh7k8UBz6wCHXzxpSxQ628YmxC/qlb84UZuqvO5xi8mtaQM7UqmI
kLGxvfmjfmfocLq+cVlSsM3iAHctj5lw06UIwCcfZvKqv/aoh+kL3S5IJh0yPRuz
kuYlCmw/R+rxPKAZ7Fm6HF41Wlzlqp+3TFWGgMwBrk1ud53VGNMIg+NBj06ctqal
CePMz4cJ54O9E8vQjdmoQRGWcIDwQ5AK6h/wbA6p2DckWJMdkkwxLo+1VfWODdl6
yhtNCcUdVmWFfd1pXQtcqwX96lp0CxrrD/Bjf0gSbcq4Qhf+R91GZT8KrB4zW9xD
Hs5dgDs4EKuu3Y8L/0dqfzkjA4jfGX7Dqk9vMAMMsfa68l3VrybEcMC4A66T7AtC
DUiFv3TJIYltFH9d6XYfWe/2ZApTE77FSiuc/0VTSvGemRhF+0bMbl65QRw9D8Fn
VEydivNsBpDOjuqua6FTtU2zGsOSLfYSKQe2h9UU/w2YQLs9plrDfHHmEU0mv4+m
nOMtSn+AEeiFul5PKGkKaQZPZ07AT5/yKNrb8Vvr01XAnyamtjYx36/TaA6xDvao
8pzAGQVctmxGPRswRmP5IgpU2JKvEXcFr0helJ7eK5zxBHCBT0ylV8OqCKCzF20K
uxlyfYFFtwx1JxHc2WAEEh6jTIdQZzDH3Cl6NIXRJwQBS7w64IpEVxaA1sSe/1nC
z9Tp8i4reUEvu7PAl7svk9a7jTqhlVNnnrRE5y9UMzQxyfjn/lfnLxcJ1lpIk4hh
N/xxCzJgisNf2pbqeMRook6yCHLlECGS0RlBTrMUDGUS0QbV0r6mnjU4F7nr/uZZ
E2TWdiOgF4+79F8kaCfTSGUc5bQxJEkEn6JFFJGnkdaa0U68CvPDI22ru2ZDkt6Q
1VqhY3gbttoFPtTbSAfYb3SvMZZZNDk1kOk75rCL92LoCF1CpmJcyDvITwd7Lh/A
Cg5bOMmza+LrBGGah5yDZL3jZkmnRNuZTHyE3ayP18PVM3H8r5nCuaj71i6zq5H9
+/07uuVhB9mA4VW7dQNj+G35HHyC7YBT05cwd+KCAMOSgsIUtECog9mTMEeXKWpM
7F+bXsQ9hdNRMO9TiorYpw4VMXT3gq6KcH0w3fNTEPI0mlMqn+UptoSqYcHOHZfo
P8sCQZRS2Q+qQ4QSkS57uf6YRiz2NrVgNMsDdXxa9xFYFcracCvdTjmTMzcDmW2K
iC+FgrlvabzJWuHOfkSlSpjPt84Zffz0JStqtMqD9Qi3v1mHcqfQ0HvSzvIR9Hni
2ytL3tZibBQtpN1gGQolNeC4FkyWHa4hQERdsYlNf6gGZbksnPHSCXgTZAH4Yx5/
xM5qUfa5XqVIxFZh03Pcr6pTwrisZ3iKG6R874ZDtynHq4QifliR5pszITvJPbpr
QtXj8cg1gnOV3T7ybd9p66QI/enawqB0GPNyHpGApzblQlqXHUsFeCDWzbQbjvy7
Le8baIlchK83OqthHuQ5u5YMB+mbfBNed6Hk5x0BHR6GOVq7UB9UwkRY3OU2rHyd
+MRpyVYGLRRljZqOURiJFo8tGMa4EpJ2udb3ej42SWunwKAKm7h9r8+8Fmb8+7Hh
3DX1xg8+XLoETOWPVSs7twMFDspKzUAKyVR80OeHJKntZ2tL/qKXlgxUsjakdYuI
LCKem1z6yJ1pWqdt3MAxszG/QgRWJ4xyTzVjPRsbtzdw4df3F3ydLoqb28wjcJgY
1rZ4HgroSdmIY8074c+34idTVIfWXfLuQiIfpTy7B4MnA+/IPTYhtSEZAzsAgogO
MrZqGVo7LFg8xe4htg/6m/mXSu7V8PAqJ2vXeeWRMeuRMHaRiAMOXaLbukdGRV8B
Zik4v+wNxl4P2JQezFUna5P+EVtoyN0rTSXy3WqCCoKwYm+80viURYwdCuwjY5Vg
oAie3HZvsGcyhYzv4S72/wliI0JmIBBMv8T3xE4iTzIWks/tHRtMB8oowO7gPGb6
eyLTlzw0fP3kb/14Igzgx87ptHnPCpzZWP0Pc1ywKkO6aa/VaZL2IQ3IsUpYr26i
DzYZ4OY4SN+Gq2y0kISlWiu8WYSv4sUUO8oBcpUpod/cvjYYLm+17PjWVI84uphM
ZzazUFYkFulETnRGmo1zhQLTsHfSiBT36tJG2oyDyQF+66ThwU7rmxjehLWpAM7L
XOnXVfIX+BlIB9kcNKzYa71q6blbRcirkQ6gakk+MhVuuL6JjafpQW7cCO9dV4I2
PhAKN26QsnQUbiM3Fy5FqEULpzVoifvo6zRohXQEkcjnfYp8Jmom8OQ7gxDkd8+M
UjxWn/a1yGXV36qTOe6EMaLm5mwHp9/HkfnUiQEwh4bDdF9zeGv4PomRXqBMf8ex
6Ud8ZYjEcvFOAXS+1s3uvgLxKb1uvCaBvGbuRwa8lOolN528kDV2rlBfUOHrNlFh
R6iZwB+pO0r46YIgY3/5bpEn42HxeKikwIJ/sLOmKFrYVVFyofhG1qzakO50u1dR
1cnFAcdJd1i/SkfQxgAkNojQIIyPrhK/WROaZFUOKZkvmoLmHGf006q7kBhfAffj
ytkcuNlyQ8/BoIQFyXCFROoWyXzqq8b8q6hsETijsbUHGaTfBKc7n1PX6YUYTGCB
xTtiJVm0imoEJWDjqOphFMrrREY8xoWpjkE3FpmltxiP2y1SH9TZWdxSh0DVcl4Q
k7c3lmX8SiPHQvQ9ZsIvpHxUH+/Z35SF7bSHwVPI2bykBhWDf80vfSPjXgFJdbE2
YOQRwq0wRbOXCCgqmWJ9MWftP814zbvV7vS5JU9yiGgpGK1W+L74rHsTIvRlMYsg
hzIaO3tFGvo1rD169VnjuZvSCJlBWXQReqlGgGmy8OWn0K9j08oGDIK/JJBKsZ2m
X8O0tqAR1OuNS7YOheCzJTx8aaf0NcHamt4OPxuFmM2hx4mgKfOaw6vfKuhCCEJb
CE1wIAxnM8Ctisoxioswb1to76A5mZvra2aahSuuWHd2hNxJlGKGmd+RbFNKVq8M
w4rvK9wHd7jYou2b8jtCWcehZSDKzT7xBuvETGt8hBLYdktKT7qnMMya5Iv8gAzY
hwiFcgBH/4Xhm3vNTvvyumD13SaIAhUZyPf7QsSDhcJL+QhaZe+8Xk/fCrsJZME1
OXOpLd8mFN3ZB32dQ76OciKkqY6aTZBSwOexraYMSjR2026wD7xLZ7+IQ+Ilrhi6
D0RsFsjuX+31ltxbMyxxAIZRYB2cHsQCQnik8E2XTDr3mz5y0wKqe4giORQsSd4Z
bj7CI2JZkMXkCXieOOsEA68XJpsbMgR9ndP0cwLDnyeR29M0oEKzZzayLroAVHp1
TXY8T+Nct3ZZgPNpRmgflQ/ZxiLuDTI6Z8dUfzyNWBzmwfC0UxOViaGt3tfcUw5A
YlxQtdZX5GHxUetCcdjjRIvIqhXJJC6xbpoYruCBIIX0EYe5V78Uwugqn0o+XjZe
mDc4r4q541reET/oT3uzRYJe/PpCD0JdSC3JrYalEtvRS65VMOREvdjXK2fCmbZO
Ig2aFN7QZnRae6gApI9XLOc0IE4hb5lTQdvafHb+yKfuj0PnyUQyg2v+W0B7UrN2
+H75JJVCrTXQq4P1KgFvCsJxJGL9WNItxJalH421GDKExLjaFF23dnUWl+lAx7PG
e7MzPPXHPXiEaRfo5q6tq0ih7wFUIZLtnO9g9FfKKHOnC7G0jbdsRFZXgBLj1VuV
JF4lngokr4nfj0ztRtJAO0x4f1NOvEHNsczWMQeyHjHD1fBKaPi7K10d5bYQolF1
otJpwsfzcq5HacWzdwRSh/2EyapoEUlVlRrQ9sIVkWF8C6eAhuMeOipSV29IS9X8
s+2XSQB6bhPDTtx7kCybWQLJ8d8T/JqCMIngWIDpT9asun7N9c5UMJwUGXsDwkFX
tYrpJo8Wts+QEC3LelTtPWy9Q8jtK1/yX1DIke680sP+pbDw51+cFjgzfpyRdGys
UdIpTotChQAoGokwedE1BxImrnrDtIWYrkiM/MkYqla+Cmmx05CDE8tDnBB6RcbG
eKHHF9dYvNdBk9MIlA3cnd6mfkH4lSaD/69RpC+tXSNhQieRczsg7Xebna0OJWXF
pMLLHNie/SNVmIsGhuPbkfR4anXmfU6g15CGW30xECdMh+hCDIiRi9bygV5goN+/
C1431HxK0xPFGBJj2AcWwaDHOS/QTmIYdhxNGcFypQ1f7ZT+LwsLJzC0ZXa1jM8g
HrsJeCnGOeS5fhtUk+R1HAcsDJOTxejEHrTCQTxdKjFUhF9Cn9feSpECtZYW+vWu
4ai20iKF+NYMY9JfFWkeBp3T6ndqRkO/Q6VyPGMiyyb7WhzftVHdpqh2ITqImWRo
8tpIh93S7VEnIE4NwKIkZJr90XQggQjaLfwmRnXTKr5nTi2TD4yr2NdImQF8UqDM
K36Vhl7kaybFDLO9aaYmj1oD5GMjs6ylKr7T33SXxvqFscxU4JL/4DOyB5wg4fDP
cF5hBFF3NTEliwoJan61UVbzt/lHytt0dxyrC5Uu5X6dbhNyqS3VIUWZPIgY2Ls7
OIacTLKABdh5EY4hmabuiuTIoG3aNNUN9hSybHMo3IOZ35sbBft1emz+W0xkfEqN
m0vrY5zJvVskcbeKaqiI4x/vMPMvwqD+o5WhQVTlkVWiA64fQHs0fbGA78W0wAA0
ZrJ5KoeMlC+bR05tIpNTJ61bo0t4/NdqlCw0h79qzOZih7RW+lK8ZE90WRJC2W/O
UpdzxqQzzbUbtIwgmLjlulCsOqfok0DgmwlNcVfut9V7PaWsc9IzAgG5vc22vYC8
YrBtrEL0MkcHnYsPcd+opb/0gSicrWV9NjpEdgoWbnYFkfkpc7aIGDwVCwsVUC85
0RXhmI92iDVw7StvysPmiDpJnGHgyE6vZxlKSDIHuYn1KwrVZFMJu39HJPxFStl2
Xr2z/AHm2xEM3cRg/Y86wesmYPpK4ad4eGz4ALztt3wyYd8xDLb6YROp0/RtoE8S
h3xiZICjeB0xeb/BTcK5h8cvQudjrJ3CPpBia4maIvjvwhRgUOY+pIkV2A6dNTBx
Vb3qOBVu7QLj1CndWaJyjzJKaALOEQCyuYqIqb8A21JUE0nF5KMTdqiNjgw7s9kr
jp5AfvSscQOwAF2cnr+qWYtYkJ3mAVAxiKHFTTG+csUNWtteums561Wc1EKSl9AF
3L/T4YdIz6AuMBc+kEJsL7PxrK2Y1ZaveMEuFZqOtylaKjH2L/UIzWks/wheEDPY
an8ygA8yp0YcM8CPF6VeAE9VE9LO+N+fmNz0FSjjrCKyEAmJ3btSe/TCArWT2n9c
Xtilal5XPJXLdSZpmKZaSpKLhddDuB21mxpHfcJ1UFwV2bgpmeB8DmkDhi4pW4Ew
3UwaF9O681CjVZQCdhZGhNck1FBEunb8yRgYad+mqKMASZP04TbdaGizdqPflsDn
B0rYdibQbbaG8orN1NOlQhIhVmln3g+NjQ/5pU7q3sEb3jfP5KRPeabFBhW4Pk1B
WkCIvRqR4ECm8bdY0TYY+9i6fnbHA6jg1EUrSNRfJL65L8HJHKXI+AnSCcucNKbO
q1cc+uYFX2VyHhsJPIQ3Bv9nwUIo8Y7T5bpH2RtLJVJJ65ebsUE6XF3a0/aohLT6
a3EMsSPWXPc0J1mxDaZCqJEJAiHfMswjfOz4YLUs4HTV6qM0d/PfQzclChlDps+v
xlyOS/HghzECT+ansZu3Apf/GbVkKQtw3d1TyYqFk3xMxGclsTKTHjMdHMm2iQ1i
yFtG5RCm9R2yeBktgpQjTFX18gx4pFALj8y0aTVJwhpBjnLPaNGm6pmUss+b9GYP
zVVAjIYhi+0mr361ACTlMFsnxnd3dmiBmZ6C6aDjrfhY50WLgFZI0XKkn+F33yWY
0RfO+NsrUiDjTmatL4+pQAdY3WF9Xk+Qmzc42rJ75Gnsm31PVmi7W3sNCAqsm2aP
ENG+ZVcRPmXJZTQmW1QD5jux58GInxvrAwhy+e0li/18Z7vsz0VHAs9a2yyFBjkO
Jc9DqdY99TYXfkHFovMEtK5znD5ackBrtro24LmydPopHzpSNTdgLAGhIiu7phCb
JMOmncKy1u/FzNAL/4Nfs49a1OcoUaTYl1099TrvatIye2c5S14wdX0hXh+DnD4W
Q1MKPGmbh2bzz5LCg9IN6NYaZ2soOaBHBdpaI2n6tD6WdABtZOfeGwip/NvFEdx+
9kFCf7RLG6szYLhfFD5fXx6ByEWAmmnUijmC9WFNd/l8ef2LFilQFJoehAEtBKzD
mjx1SiY3rhu/ct469OiFFX7V4/mHlndY/qCuo8ETg+A347czDvjo4g30DXW4yPxu
iYChsnJTOKQ1rctSyY3xQ2BJKw3Ci7UWOzlldEsmgHdPcL+hAKvTb9vrqMx7lug2
ePUKbNGxeuWjIDqMzA4vBHrs0dYieEwKDd//Q3BSVzaZUAXY3PPEagiaZ+CWNNK7
xsbhWYwUUxHN+aEt+ESSTT8I1RDcksf6ixpYPUjS4tZ6VZRKmh4JqoAs/hN1y8EA
e35hTU7G59Jli7ESE94ZTWr10gl6TN5Bkfoe0R/iEB0W7CgkRKYDNSyKnnP2OsBf
ZGhPG2h8TqJQ0cxpwoymJA1NRyu4vOllTW6t5WWSMWEKPENgLwma+ug99WLEjozG
zu4BupMALPtivXifHcW5H4SosUC/jUZ9okMTAsapQ2KS01g0tcP/Jmo3FkAJ+vQN
hqn+crwa4FvinSPYGTP+Wv35QFe38dBRzF4+5kwfwnCtV0hbYV7cKkL9R19JOWA6
Fu0POp/HJS2QkcfRxqxgFnaxGQs5Qw2fX1dsu02HY024zjscQSn+13j/c9OvXgee
t1/IXhtfnm2yIgSulRpvu/l8KgUwdBgOAJFuRDTSSwnEOUWMgW9zDyFxPcR62w6X
AeQq9mPeHr7N5vsMh4UTX7hPj0RuNGI88ol1n2PTqz4bqW+sbBE2WWWJWxHxt5pq
s9EtE8KSge1tWLgzWkLh+DtASMqc2YApfpLrXFsMmcfvP8m8qBbRGKzN5TKP8O7b
pfPBg132JuD2W0oXNmGsgYDq/W7ItoyxYT8jzrFL05c3+C6CGv2qGZpbspNz9A/j
Tuvp+U+3xWhK1bKp6H6cJd8b+vkLxXQgPr4DNDLEL/DXFz1ki1ifcRlfXsEO0Gsy
aKOf97WbnaPrsAgSaOd/Uk1CuTTCIjoO8+SvqdbJAnNb9Ig/p7wTR2vneOKCUfdD
OaAlS+Z3YJAJ5S/mLBSX1ySmdj7OvJqiUg+ov8yFVUsvAKL5sCaZWgUuF6Pzgso0
vyAxaFrr0VDoV28yT91lnzvHQtUP7NG0jihTIz3A+yGqnnYdRWrFMayxtIggzA0D
suZVzveIr254bK++GK9KjA==
`protect end_protected