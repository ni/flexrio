`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3824 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
YachDS4bpHRDzLXFQC4CtfRhLaGgZ3nLRqULRDrFUaM1QNB16Zqica2Ky1bQv+Gm
l/3C6W2voOoV5VByJqvrSvwwJk3uMRTYBvaBDF0TeMGA+1GKBZIPbrpbeA6Hsr5R
MGKvqvc22W2sXJoCD/UqEb26jb5t/YDmWaVtwuMWnf+LNhlQnQa2y2UGcRXzPTTS
VlkZn/D1QY/d8FkByiUJlstm7GXj+WuyUsSgFK3HSccfbFrnJi9yVq0BlKFbgFGl
I+s7YPMz3e5rZW1Foqs/kSpVHyMyZW6s/WOav2dSIbelXFjn1LH/URRjUSk9G8ZE
vQXI5eEcAvWzGEAm3EixavsmUMXLMd9cZ/VdWtksL2NIxdcZp9Z+w5D5Ie4h9ryN
EMMhScZ9Yxn/NdbVT+sa1ql3qCJPuyMPDalEzQHXTXWUbtzRP3X1xfyHAVgJO0CX
Y6Hs5vkTGqzbRp3MlqiRwP+xL/IqdvQZVwx4XsgiO+pV8OZpt+KS1hU/WZhJVf4f
0FoGfh8rW/Q/MgQfzZ/nJS3Vl8F8Oc5R6QPpHc1AKeVWjThbMD2oHPchlnyFQpU0
E68QyHrkHrXrZKi9OmquznauE1vuCcEqda0sE2QuWoC/rj+uwf/a8Q1D8aN/Z1O+
J3xiOBH5zdj0NJqAmGTxEdo7hFejUJjHhrEidjEYeoVpB4plMj8LKpM9jwC2up0R
b2CAqlP7kCBwwz3R/Zny2JkJ7ireGxO8Skgn75hd3RW2pM0b7kmzghorfJ/TLBzD
seklmu2IRnCrRTzyJR6u3d3KjXx+Rne03HY9zE8ieb3DWTZkXjMkV2BiFc/7QeRp
GjzA+g6R6AMHci60ixtLEKblYQJ417jcVm7pwz64Pfb5soNYPhZkJ60GC5+xDezQ
Dje4q9pzZOwSgsAOZt2iLAH3gFnfKZa5f4IU/L4Aw1H34gCo05CYjx3ZscTotDWz
ze2M6TnpLhS8EWK5lJ1LHRRViC5ymHT4Dc27H/10k3EVvJu/GrHz7bH6fm4+pcvg
sBZY3ohlAeaivcbsNpiw/151RhJmMdgtUuqWUhsfG4vw3OihDOnkWPllIJeXDSlW
XZBAENn4mgG4aDxuuS6IVM7c1gaPELJTjgjcaEGccPTQ6oQYrOk4cOQYU9hVzH75
CaSsRozAJ+D9WeKCr0bQgOoT7gSJtCnSMCCd+N7Wre9yiGZASMwIcBsHVbPMMHVv
MT87s5UQbgmx8sladgjHAtbUiF3fpJFPxzbnRaYtNp9x6dLuPOIEMs6a0MhJawxb
/CGf1sCQLIWsEOUd47K8eTkMNNAVw2LqfPzXi4jpDDYbn//uifX271XynjhcKFqg
DXBRMKGFUHLbrU8lQDqAFAzoO1RGoAaCZKa5eb6cicxza4tM5uljnmUrmtXSxGAE
/PfXNSlfCUtqCbRNKYkWibGJvnt84GbU1pJyQ1uM8nxraQhPzvykBUB/tcjt0PGv
3hhZCDiKhERNlAYQc5xpO/oGUXT3V0UGm9h1+e4QJvotZ1m8Pjr+EHuPftNF11gS
oJBa307xk40WuFf4rVQ7BCyspzcDgleDXzCOG8fln2Ak1ZPraV10M94j/uoKbhg0
bQM5fJilmeHpSwCJJLAuKdRZBE5Ub84QaOZpd5I4R7WQBGfvsQEhb1OBB+b3XOOl
/fyWY+uxZgPXRjSeEV+JqekCP/mNJI6hrDjkLHduGuYQwVUFN3ygzvR+XbpMueJW
kK0MOVp3VmH4z2PAhVKGup+bwDiqXLUM26Wqcrgn4dnu2ULlXdPXyEdLcftZpBBQ
/Av0chyeY9E99ZpHHq6wP6phu5bjVDh6GxjuosFFHw+u+HbGzbhZspOeKo4bjyzy
rjE+ToBphqlFobNG/GYCgFVMxRFCXx3ruwdGRrVsus70gaSV72l+vrHfxxhYH67b
URjgMzhGOb94vxhQBze8rX7QihJVy+VWSBeY6TnQLdpqNBteiE9ZGwfaFXL+c0/P
cUXATzBSJb3NpRhCAXS5Ue9TISqOczG1Dv82CeFVAX5FoWdsOANe+pEIlrNpg22k
/sKXl3dr58SjgtMCzDYOF4jXt+7QzSHRu+9UgMAXP8IxqTAUc/llXoU67479mRPl
Q5Xh1AzCbCc9b/ppz78oZYjUb8YAQDcgpDjxk0jv42n+N3tfRM/IsGmPDOeayyfW
ILJMPhws9xfqzZkc379nxK9VUOEyF1G63m31RhRDvcaAkfnDHgsUHsth3P2Py8HP
OFtglVOxzmOFH3X96utK4qLkoQgqbECoXR2t0sGgItVKawqYvPAOByLQBDoMJT5F
FAuhUFNy+JkBuF6n22g3V0+2afj9puPul42MGpuJcsMTKAtOHfJ++GYDItsHhTDD
/jmKhOWCHl1C25g/lj8zJVNEVI6yPtSZ56FhTSyg6R/nPMFSs00cIErNBWRfICd0
MLe9Viiy/aUmNo4rJ0W09tsIZcWz2vo2FNTddXHwIb/4X5uE5SO05dzS7bYz/mOb
111itcbq9X4tIs6/IuZjE0/Kbf4x1ZZ8q0eJcJfrF6XZfbp1VUenhuudL6nHoCVp
RTLhVeW2UG+YSk8R0lfRNia0w4LIugcwOjZ2PALP/kVZDQXXcfwwacQJkb4GF8d7
toLTQ1N1DCTWSEUSiQB+RwlIoUrPfm4owdF54OM0EUKcyoa4nZ+4IQDUmdN2zdhq
rul4FFgsSNSU4icCVbF1KtKjpGbqDjBypjbm/KV4W5S6qZIxcSXiytT/lwjYqdyu
PmeSlfhwwvPrsFkSWhhmR/bsvWEeLidRYMP2tUQjDkw7hfzBTvBmdt0zU2T8TWJz
zU2jstkDJRB+w5LcwZhSB5wlbDuz+xe+3n8fleAnNGmM+bTXikfRoH1HgbzMqaaV
fMRSykpb2j4fJWhNP0/vDK6BN5U/lzzp3jo71os3Y5n4gwa/yensKvvn8kvLtWPg
gpYHlWhi8EYYq8YPvjGkBIo9D1GZ1om2dwzfD12bghicOpL4TnfiRQZ6IvH1vPtc
W8VFyEesZ8X6BteeFgt4r/hNb0gmX4hEZwIaDjhvKwOyTCRD2kDVqvADKS9wM/9e
IFgD/Mo5oV30AJMnYh+/Fvk7uM23VXrpYTXy1TO+lTMUDADBhctIQHhSnNvDbSeW
jEdYSm7ikMpcU7jxKHhFD9htJEuyayMNpowhCpWPeWvmjUVEK3OUutf0q5x39cMg
sTQ+RGdmHEdTdEWrlOxuFNdGaMlbsAkCaVKCafiDukc6V47zSHgr/pxXnA4S8LIM
LjE7BGy/ckpizVc12zFr4riDsozSu0zTK4gTj58xuQ+1j+Qukvj89e/l7PuP8TiQ
Q60htOhjMr3WQ6CCvnHY6LPKJKhWKol7JPWzvrmWCzjCnD75KEIuVdUkEyPsiBEa
+cvjXk1yMtxvm19h1FIq8LGMfrYejuRjS6hL2/p/steNNJrxY0PWTy+zi4Ioon0v
kZo40DGgpVmiUSQXgIhwWkD8PaKJPRm4cxTxQHjOMPIkFwDYXjqNzMYkMM7pdx5y
4wSp3v+R2IWC3gD9p7mpzQdzJphhB2qQ/FHiyj8V7Y9Nq5eloESUzR1egxn+Sdy/
Mx05SgRGCKtr8IGnYWo1cIHYcnTXscKtebM8gd5bO0cvtfa1E63lUjzLPlI9jjgS
Ybs1O1UCKdIlVO/f+fm7d66ofi1/d8fR/MtMYWUE/zQ8vx8C/R58tWhFnsPAwlS8
uqSFitfXO4aa9Nj+6ywyRffrkuNJ8lYX9bT+urHJgdOLJS9p9O5FQKzkRk7pVKUo
KcYfViocwFkm4nECpUaoKPWkoqTlu1OL5Zi6wgPL3ThBrMAm/G38bCeruI+3LFkZ
k5lFBIQ6dFRHhBEUaqz6ZxMJeyY2OP3q+0GtjB/b6VLBjc+h8NG+Sgjm7sidepzX
7RmqjvTffEa4ofzg954Y921Lcz/hu0oec9BDjlktNX4CieHfvV4dXAIBIB0JGDuU
Jz7PPRy+xX++Va//QsmjVaxSy4epv13dhVbIiChCgiexCWCJlC8pp8FpO0o8lyzk
XNDtATlog1D2qdFJDUL3iR/zAar8CDd5q3qaxGQ0FB7jBCvAfIGEk9OpLQzM+8RY
Wsu3AGsAldLH6W1Dimwz8gB4ilCI9L+foo7TF7LiNiS2BQin/1f4PDhi8jCQb4NS
YTIvgBc98kbVSz2wrYBPePmZPNVSZOYi7fGEobiyYbTwblrff9WChpwN12XInrnv
5Vw+o5A+FILJKO4AA5z189z09u5WOSZUnOfhajLvv3Q05KHpWoiM4YQTlMvlAUeV
j1eS0EvLQOD3jYl0DpomWlzMlgPrUcmIa/fOGDEWirk4wvxGPd/811mWvXoZXmZ8
44mOQVWbGRv2eN6x9bIuyMY7QuXF/pnrjwvYzftMwK8lqqK3kK8iukIJYSqDI+lN
QsJ4aF3+ce5CMhkBQrzg/VNLCrAbSF81zcDkz76ACE/HPqKH7zG7CvzlpOvTJME/
uPXa7SW4vqY8DNTF8cX7ymXZNZ5BUUJ6uf3DY3mEvNEI2dIvUt5oKdFctjXnJ4qk
Ok1wJgwEgoqrygeCUS0p2zgqM6v32hasR4HCrLXHyQNXLIe356esFnIWjr8ZBaMk
yeNN8wPNiwa6yPfHGLrJZFR+h6NWJvHWKvllUo5tLGbvvpI9rvsO+XZeQuUT1x3G
yCIXHUE/88M3hDG0uXueY5Bm2PF3vpzC/xEMlf39LaATyqz1l8l4HZwarONHi/u8
kks4rVH7Pdgmx1MMonR5GqbpgGsSwS861KZikY5sdIIN7g2DWwm2pmoAYAIJyhRQ
xwei7tn048qjEiKUKThtHqzwDfeqiodvL0G8cH26KB4kWZLHgnlEmBj4Aau5Lols
+pt1Fj0RBI3J0H9a519s7dcBl4RLN4q1ya0E1CzgUAvLaz5mlcJsMRAroSfLuqPj
i3ymjQMdgvbtO4y8122Efa1uwLYqM2KfMvfqJzV+Zlc=
`protect end_protected