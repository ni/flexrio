`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
dYVY1GBMsK1ODCn3ZUp8SoAWP8Fvt20jOclKciHf7Ysn2OlvHpNHbXI7BFbSBeZ8
c0HSNxtSIQSCmTTcVbiOe5bNYdnShY74EmVDlUagwaODhK9Urx30VHPfg7K0Q8Dj
u4EuL8LzGtWyNpPuuYUPfH/EWWJz8j2B3GlAugKl7fR1RciktYEXyNArDzj2i2Lo
icoQhkynNgC7v9DkMLR1BxAwtrFrckccZalCrbzlnjwD/DOLPtfjLaczesJPkKoa
xZJUnnMJHmZHdGCWDxS1eicDF7kXXzsE1BA2jAX7HQtg/mw+vmEQXKqvkKy9tRtW
yhUEHOXSIVFkC6gJ+buK9Q==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="SgR4h9hEc61j3UcDg7JP89NUc7gPf41F4aolx7zbZ/Y="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
PcTZf+e633x3tw5Pd+98Hvg8K8pEx1TP/UFyHup9OvIvZyp7VdJ/eQ7Czw0TCb/d
NGL0fQmqipTyP1VBR/CwCDPv8pUq9mWdoIhPzGBVMq1ZfAiLygNMWUwFu0/xPfyw
rAKvJfKF1tLDCsja4oREz1+w00FDmJ2gsQcbY/9d4Lw=
`protect rights_digest_method = "sha256"
`protect end_toolblock="fB5pBzxyhRsqq3gFtq6qZ5Drx26WwP+GzJuJsgJq2oo="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 38064 )
`protect data_block
Pw0LuTSwA3gmWF21w7rVYBcj97hqvAcf4dxm1w8M8xOO9V5Zp53fD6281Uk66by2
V+2le3pjRQ4JkfVvu0vvltrqFdWvBln4SM9xPIyOvOjskVz8MBZo3CILQk+Kjz/X
fnbKbjecJcaTOqZL38FoHcql9OjzxXcbVO3KApWzB3rFG05wQmjZe2NeobDOTDFH
jwqAAqIqMYZ/t5sNsDSHFog1GzmuhsPvqc8ObOUzAaHJ7zl63l7vNYSKL7FNZc1x
2X9IKuhCZLuT8iNCij2ZFApIBOFq6pZZ0LqIfNKJ5yOok+tIApuB0EKzva6Xktcq
jBjSQ21OMozqnaBxJHeG4PWbn9m0rsNGYN2rz2JpTWIX0dwpez8KBLVcpulW476f
kPxTMr+6S8+Dj5SGQviyDtzXpAg5CkHlxUPLfPwwnnJVUnMC7Y6Q97r3eq3H4G13
YXRtMA7SkdK1szVViSSx6a8UEjCgJqNBELys6R1HCZSZHnM5CcVD288u17ZGmt2v
7le9Kdr0+J56AvhmhaTho68ZKp/nd3KyjjM7XrZCDcZjMkV/JFxtjj15mOqSu6KU
/8xlxYWBUINqYBn/E4BcRH6IJdw0ahP8YatdlY1T5oWmotv5UMOKwTScyRCKjDd8
vy4cabbDgE/DCWUyYRAU5K/uGHk0+BkNnEb8FTlCJ8D1mGFof/DOYr0sxxRkA2RI
m4JyPhuHAdc5j8I43EU94zcYRKsW7zl3VTEk4Ksut18JU4CnhkOFGCwwIClY+14A
GyCiFMcpc90NJJmZxkUD7q5NdEuirQbkH+xc+Q5B581Vo7LC6+z78JpsY/NtJW6c
OwqFctjbxEJrJZLTXeEq8UJk0xtAJoCzynu76QEck/FMPBJHxx+a8ieCMEnjLiPa
RPwQPdjyPk80Q3XXsq80FybK8tg7U5YdMo0fChno5RNLtz+BW2o35KvvMHfuR5EF
zBg9MpRIpXOd+1m20D1xCiAi6JojdIEsMw07ED8wDcEZPzveM9TC1uSYfeSzrb9p
HTLxtpf1oI6gEZ1BFMwujCSXfqone6QIc13tQfHNXe+O41F0NpHQx+6Ra5WrgE7+
ppvNPUDkfL1KuBfnYiZ4GO46+TU1J2XBHv453inWQqB0OeatS65CldEedEbj4ITn
D3C3rioN8yWzMHvgh1VW08DmIffUYYbTrBpGVjBROfwzHcrxxA7f6HkvOxz5u6Ha
TKO7OpqcPm2/9pJk8l/o/MdAmfRn4anL7FyRF5y1dznumH+joBKqxL+VQfQWpCi1
xYot4JGdtr2wcCzCqWbUJOglHQmc414jgJ4tQ/GTtztt78G07+mwTXCr5d/GPegE
WARXsMjrNEDpZRLckScuUblZuOL5OK+J/qrq6BppYwhq3OlUc3G4eVxCW5oK59B2
iIy4+3XY7bF6+UPdizyzEf/0rCObUqLMTn3pDAisWOM7dgWUPgfd6XLk2Mf2JF+m
niCmysO4ZfrIUqHknZwHdjUHSCR0zAB5VU8xmxNq84i0N17qwiB6oX/lzlVJg9nx
5SdDRfB5rl/vWu8SBQ4++xsIqAHNUWtg8Bnwa57kBY1sUvI63Exvv/oSIyQv6Bgf
ovkqXrqc7F6IgVterMi9hbW4hXL799vdyAdQ9giZSR2xOSx/VmwdQOZTMtvkZcFS
dl7WYPxmsv02ps70gnZh5gkHcDBZXw3gq+WwxFdswh0hyiIGs83MrR6pe9OdabBg
dI4uGudoyCx85YOuI+tHyNA5tIxQ1qKYanqCRpUzqdHqdV7RnNhEwzIIVYAsItK9
YegvqbGs/a2NQBCnITv0M2Tlb3j0cT99+9wdEAfyhPc9HOVMAx4fdOHYxcW35g2o
DyUzEe1ZQv0CCrY6Ye0+FJ3iLehe++jZnF6aUBG8Qz3RHpfUyZByEDRG1U635Uf3
R7PcKSU6jmD01agbo5qgK05l5MCgV/eyXHpW+FiYyozpfIM8XXxUzumpaxBVyn2n
tGHAu+IDcTG9FdXyXxwEl8caFWGisg2DW7WSy4n/Up99y5G5rDHLTypOJJJxSZye
s+C/FdBpby+uc7FPGEX4MCptcrjdLN/iAka8sZ0Va8oolWKwSBUvVZrL15d9hgHm
G+tc9Qp9kuqysXAdO2+6e6D+ixnmfaQm3WSaYQ5V37wX0L45jTfdoQMQyZ/9oBBs
q2g2CXMImukC0gptBAcpHYzbt7lhSfJ64qnCeXo4Q/VkXoCbSQY31jOCleLQu95i
YSVrw7GM++Av5Bnb61LlZmmaUJsFe9e7j4y9UL73b8urPh4HAtTwg2IJZSX2tyti
bHulZTsvaj92EtvDxStTSIgFq0fK33G3unHc525TUcIc1D5B7wACMFVYIcfDXAut
+8QKghOrvlP0hFYk5z1dhN/DfI/pOq5tPgq6Msbq7Y6jCtdbnWh95Qt9yn1t1mPB
9vDqrB0VOLkA7bDtCH/UGeZRx9FFRK5xsStnzcQsHlRYXF8uV+fq/uV6uzNQvct2
HMkXRPCqReHyoeUxvh8HIQglysoOU0JarCte0ZStuKsJsyYcRIsBfdjlh8IWYTJu
GyJF34SJ/IOQrEwnNpqwrDMa12JIU+wK0yFmsJFzlXEox8WMlp9qclwzioyTEF+N
vb/NV3DsaYLJWLEJLJb0aQu1po3PfPZcFWnGPhasfypR9z+jSWpcYcMDi2//gZJm
ur8gaMSHM0cQ79nHVZhRl+jJEtof8Ahz2fu9rYc+E2uC0Q6LhyG2+e10G3UnI/EN
wwaR60fB3zT7Qj8+jX819oDqFnVVCeSBAGMbjiTaweqBiMA3HjD0RZxXcrM3pzRS
3tABX7+RZA1/pBv0/J4HMyPkm1/LKImtmIzhBO20BMxChgEnMq7Wr4hGVobuMvvr
XsGyOlUp+bX2673UVLcEetwa+oc2Kitwr+7YTp0U+rj/OLh2unF2hLHukPQyZpoF
gE1e/GHRetwxcq34FF09oUJzoRB6saeFw673YG24cALZ6h2qq6O5gKwUkbuA4lWs
JlhxCTejumoqn3W8wodYQoqu9bIWFzKJRh0EOhkBvkYACJLXEe4tu9K1U4lNh3PW
HSRxRrnhrjeo3EhBXqotEeqcPWyXFe9EPRv0Kvd0ktiUSFTUHaI3WzZva77iDqZa
lrLPJMDYUVKwXOxGGhIyu5dgCHvkMKn05how6Fw8cpbYk5XLDb38luNFNR8YFvbM
sAJI0gF+6RAFMM4xZRrvZML9gYZ1hrICCCYzCuOIy4mKonWgwSVtWM5mKKhpoUvu
xFuh/KrU71KsA+8yTiHQCe0KfQTlig/aVD6qN3RhAtTUFEqez1T6RmZupow1p9Fl
Ps2+ocqPl2xjnKjipf0QPUpIkWifkCjYaS9GMvEyGSViBZ4T/tcSRNuJ8QAjpPmm
oUZtEDINHPdSJqJ9rj35rSgOO20UbhEvS+uK0+Ls2D2/nUbpWqzqqspswBX/wyS5
rss//KxP3ewqSLhdB5uLGkyRsAf/S5X1pPdE7/+GkfnS7f7Ph13uFEkz1EFzATq4
1Vp7YO8oGu6bLB4XUHvJR5FCBV09f7wZ5d9QyZu/xbv1BjWsWaTdO49oreA8HW99
JvdDoZlbJNJ1Ay/u9wOvcIFTBgq6p5bskc0pqOnn/mDbymCI/N4+zmBtvtWIZ8P8
f5nw0L8pEPJvYG+MN+xlAaLX7VLDQIllIkfK1pYVW3gseXvN3o4yAqxYLLrDWnjI
1u66rqDGLHmWH+l0OzCjnJP8c0NLsRViUPetVa3vdfV7Ny1mzauNF2/alUGj7nNl
oY48ZROOTulWrmFMOZryE+w9X3m1Wup+5ATXxq/lC+/OG4o2otNF9ExFl6QIlGtx
BdGWJBFRWgJMzZel6vt110mYNMLBpXCmQDXLbKQwaYm3fASlzwubs+MAbUoS1N9q
947qoxdHgsmyDy10+MPfsezlwViLAjLY4SyVeJKoTChKKAR4uPKgSvqnLB2600Tj
hPg58OInIHSi3I+pWXqehsVaGkW6qwRjLdCDzwhIPQjjONtpp8IqGImzZf6SUM3z
5kYpKOh8gS0VZbSu3d/jfE9P9Yvl60lfgJ/BaT3ym3btZte2ZT4aliT8rg7RACZH
hsSw1tmIfjdsvSmWcgItVxX7S9X8S6RScL6TS5sBPZUZFJ3Qq00oQu0lH+YiUycw
vM1zuI3z6X2Olx1/v8n3Sc+p9PCSg9HCYdvbrMMoTAF0PEQUE79WUdWELmSwQopy
zb0fVzf9hyx03LWMpWR0YRgVG3ZQN3/CwvGBkYOnhC1Rua1U2vMRbOxZcyZ5B3oL
6ie8/Omn54S2wi7NiA/571OeKiNy4QWjx0hOnKX/bdHEkt745iftT21hpGj0rRC1
0jjY2QDku40WZSDkWputqzbL0dnXlMvQn2E80hVPIingLYXPfrP4GKV3hVdrbSIm
QSK81PrAW9cHUGdTW3dcYvU419jy+ItCPK6iYy9Qm/KxTCUj2whTsy4psg18tbFt
LmTZ6HTdxrSP6scsu3xQDg88peQ1ptFO762pnaN1JsmyNRUzrNppYiMFBN9aWtwa
NO+wMENGU2RYL5gcyd6YrGzP9QYXjbSfKMxxndbq3Qx7JF1j+3mhQNB4LfOykTSb
A+o7jg5ikZ/m/oLgvTlCHH65dCvnOgQRjKXnweaReKrR14amGCOq47S3ZKTEzUjn
qkLMl3dMtB+ql2iZUl9wTXO2dzQdj5kD4tucwbZenVoKVTEaoGumlH7Xh85nFn6V
RVP15lOYHOLZ9dh1Th05XjD6jHczxFytiF82uIg4pDoWFfBNfZuuk9qFm1oB5fjX
tYhw2keY3D0dt2S7BgEGGJdmkhoD1zhP2xOi72r8CtYmzQdoAba4qBbsUlIdOAW8
pQAUQ/ZUJC6jn2cMBYiz36N3aqyzKQiMvaL5rDMTsuY4n261aA++asjpwAACKGwx
6Ylre9Bu0cjm/XqH10l2wv7szyWnGVOZihJwiqRzeCrFyfZrMuPYlGl/F1onMAjW
zcEQy9h11TKeVN4Kv53CnIgeeVBqGSyxDBza9yX6H9HbRfcZYc+OYPcH9oh51t8t
lEVBcioRiymgqk+FyGgb+rbU7nuev95d4ps9V7dqdOO8hbHQJMQZoxaXkZQCze94
KIaXPFGJe2Mric2KAQa46qNfe7f/BVQAs3CFpFd8uNABqTsgLlyaOIJlgxh4pkE/
YglWqIr3q/EqLgbl/SlVBSWWjU6VFrTA1Mgbi4SRQantSmM7L7vew7cFYGD81Ruy
iYDn1q4wvIfl7YARRzTGfMkolqR5615gcMxDKZ/3TRum+Xo+jbJjOBVFqaP83ZGQ
bCmJFg5QgNwFJAwYm5A8i6M2ASmE1r99LEtVL4uvHgFaAGlkTlhhgyQN/3fUXDUR
C4AbbjwevlOkeBdo4qq0cLAEqeRN5yGpVqqIbD6CE9AuCZo7ssZn/3d6qVzXPP9I
Jgw7vRXEiUNdu4QWNGTPIs453KK/TqmYmj+ME0SpmDUrVXxQpEI/VTqjnmdHM+7p
i9hvBa7AfCk++EZH96Gqhv/5uICjxkDyO76Z7j7nbVVzx4frad1nhBsvsZVHZ1On
aQZDEz4DLe1ogR6w4FF2/o+DeGeAnXwo1Rc2KBUzzLg7ZbC55G1eNcbNEyM66inq
SLiQCgQUEmkv9FNp3UZOGyL1OWfUrb5UHS0ir3OtQJOXKLP61NLEqMAeF+Xy9zu2
K8tmo2fmhEArEx7q/o3vtzuyJrZnpD2TR8WaosRNR6O65N4P/VDVZo3emSTfCdNs
RCx7Dh8npUYKv+8rDgBSgqaylGRc09Vl/4nzBJ1f0FVTxKO/+08MzAjjamZ4KX76
8rQlDGS3X975//ca7DRrvDt8s2rw5x9P4cjpPSXu2skqIT5hia/8BbuAVIol1apr
1IX6Yrnq+436b35X7Pkk4nQGE8DVxJ+MCppezKMNVoXRw8JyThOh7h1B5NGGE/NV
TK+2EiAIAA87eatT1wcOYnxpPguf0TLycDq7VFd/lQN3Kixvo443qfmvyrghBO9v
bcvgpzgN+B+u8APabQstw8nI6ZnDbFstMYknKQLi8ET7T4iCTH/ibl9aWedgjLV4
TbQXmxtr8e01qgai7nMtTkZ4CzNp+XcD7HKDI58QSl1zpU1aTTecXdHT2V6ljmQU
0hMiqLwR3oZz4tk1nIqw5h8vODSOyZxE2DrDNNOg5FxPVFa35Ezhgrq55Gr5oYlD
rlLL2uVFNWSvdcy10HmhsoOXYBiAmq+mog0xtXSktrmQZa4x3uWmQgCErw2iMAxF
FAuQKgXgjTv9QpstmGGoN1Nxb2662TkDbBj83oiFULAL32MfTolhGbCjbd6oAzLB
2Ws84yeKOYlOPo/PQb3du3hZO2wm3F1HnD3rXOsHqJIQM696ygD+Khv3mliCSfsz
ih4rcwyPQFwNDUE/NkzQTNwkcPMGETD4ROOYF1nahqxN94HzHf1RmIjw3yWtuqu0
og+ciLyeU6eddSiJcvFs00uPhwLlGvz1piOjf2jMuCVKVqNXqMqMWm381RbLzJfF
6gFYQiwafK8olWaeAwRJ2q98f/s/JtjdYKsy0/J+OCI9/HCJ1Q3Pj4KbdSIfHql0
E7ZHWQp+qftq4KITfqVwqxHHX83N7U3GyLDgFTSclD5M07VM816eSf7Z/Z+DasEj
ZtP3py1bQUhHNH3NvAQMkjrrRX3ipq52wCSjS4+hOkFyVIoZ+LrEzQHie8kcJPDS
6leMJjAcSh5XKP4nb2YndDZTNMc0X+0m1jT0eq8Qtrpo/3Y7w/ofeXy1im8yqa01
+3KswZuS4j5Mkw8Anv6xwoyMXCowOp1qhWvVTUpKBmNmqVoe+oABPWnkFdlGR1b+
gBWxz/LeKVyjIQH7Lohvl3CNnRwxWfsniAV+oQ/L7HWvDID7FY2VMSPRNb4mLWf0
y3WMlUZJpCoqUrn23lpfOPb6lS9f5D2Jb3SYY3/ZpCzCmoiKPxWXj7pj3F3hKA2n
fNNc9Ih5KHpE0/ram+hSfR8COEl2McodtVs55OQSVr8yBKekDdVc1yL26j6NdFyR
KFI3tPWHPKlEqCazPP5vJdzd5Tffmm2sj+OhCkc587LdnP1qwFAdL6nQaVAy53F2
G13KgQl4hsAVNc5VMOmQtujOfwan1XTJnAGnQqYyfbHjIB8yYQLmk33Dfme8JmXr
nuXoYFcLxR6MLf/mKin9SVpnVZ1BQh+Qs0xAvfVKOrPfeCBoOlcHKBRg/9uBgm4r
Me6ubFPTQp8KKxP8vPbkXMCZJohEqbotXaaVi5q0zZB+lD/kQXeiLjdxmsm/X2Q7
enSddTMaOXLaLwBrqzGhDTz5nWlGI/wL4IoMgf2gtnZtQQiPmaRupB7VG6b/ivUa
2TGr5/YeNfXX6VcFan5cCcSx7yIfk9Zoc9NoEaorEMudnjnPzGSbKB3mPfHITeIu
JFhJcT8qyud5UtBXUPeF5bV8/AySQjX5U68WfwSC0fSbBALfywKxOZtYHOUkH7D8
6piS+DWAFFmjhAVsJYkHDL96iICmytFbIMC29Npr6kOTA5D9HXJxyEqyNOSn/p/U
hIk6ViIq42nIDKbY20ZiVTA/N7z04oBqod9ndcdGmhEF8+EH8pD9cuwb/XD25sUj
Z+UmWsPwHmyneY6lhgn993VMGL/yuRLBs4o+aIczSaNCdWscpXM8FAT6OSSgh88e
Mq2uj8rJBe/RIgVuQJ+g2JpWIl67wuawcogx3abhxXfbv9E0LhjJKy+xfidUXDRX
nGce2sZJNoSB2vUAI4lUqMMYrsEUCpkhXA5QMQWPsJ8h9TB0YGcyzl+WSyNtlTG9
0ErPXqtThQIYScCTmPIFMghnhbQpw080Et1705GuisbUI+QAe0hgDjp0ub5uQZVk
J6CSvKnjbwtAfsAehih1dXfKDLX6VuSNb0nMxe/2EqaqD4V+pxpvoKOvxCr/JByk
jV1ZUvIBZnm5Q6MExRPmmAUfF0d6OzZY4Kf7B5y1ytTaMosx+5oMARBXYsgPrbAE
d0nelOfoZBaFmIcdZ5vDoUgI/WeQLYQC3BVeuqfMIaLw+tTTs10nhzeAbOoQ6lHs
ShobIbH0TDwDYDFC0DOG3U3ydGGi+Ae7WEjF0S07iMvVrq3rUarNaGvn8YD+CoH3
yEvrzoeJewGJ+r0bOvXDQDuz4MfrIhmizLw9N/SYMnZXFf/Y+3ZH1MMICrCoDyPq
nWLWhnNUgs9mXzPI39im7WiQskT7SyCKtvX6AZ2oYYTMF7lRIPu82olST7N+in9h
JpbWrdqTeFhxU9TwNFl7UUD0MMXK/33yU54LVtBrYDSbmRtDhnqOItF2Z2XEtUdm
uMxWxKPNn7tYlVoyT+9qfY7ELDjSWAOnBvuBUelHXBiS70qBAP+vKUV4gYmyecFy
2X5mQvm0jpSc6T/izsgZlVYcKnB3o81dHbaH8exkOIcgSGkSwx4BtTdqLssvvJ6t
A/7eW8TJmlTggkGGGRO3duS4sNYyswdWMuxPXigC5n0xZQSuI0xzIGz+4v3hSugo
yJUpmOKlJJN8eNaj3h/JGW3UUSH5tzFzVvcm2iGScGD8/FHa9y9szWJONMVGl+Ci
lMwZrSMdw19AMwC0g74hp4vbSKlFl6MS73Sl1qClj1lGjqbpFrubzR2vG/91xjx1
DUxPiqgACT/7LaoHmzbvJ2E3SJGC5XJ4vc9N9vIgUeL8Gx1yCWmdpVX7Yg+tiHSs
3qENZUNjzxLbddvmu19Fz2gE6HxwxeiX5GeQxXsFIcft0Pmrw8wBme73lAgn2+bi
Q6xm7E/PJD6ry879brUIZpbUranlb/OAL/viEhchLyoD2WICbNpS+cWFvGQ3gL9R
jsMNJeM+wTB1VuyNj3REWSlGdf4LrSMLvSAk0cUT4llEBY4Q6Xqyu1eM9cKI8TRb
K0dSjFEr/xF8CpDjhOgJ6TKzE0oeBaj+VzA98TipMI9WUBA8bpAvUKB0ORT+JUxj
mQ4BU92iycjlRv8jaAnZPNeZb+8ntYjgA7c23W1uO4OoQAsMmrlAIyfo2Cby1iTb
xVHXr37DVKyjwsEL4FRnZFTnGgr52nLK3dw3QAK0Ah0N6S4L0ecQBwDBSxw2+ubu
xVwr6j2lyaL+akuNTalnHubaNaW4HWaW6RuBkFQ8RwZtYfKIVgSRH/ldAN3wR2/B
mUN5Rw8G9M9lhOI4QJ/RV+zdle4E2YM/dC5Et+kbVqwvUGhxNI6qLjEmeQHyeH4y
GatculEuGI8bGEmEw3AJmciYFRMDmKcqWiAsg9ZtycjrsiB6NMZD5tK+FEE/tzG6
zUovMR2c21EbJ6H46SEFv0ylb2IeyVkVvEPUkxtCegcEEP7y7E+IoxYe4zf3l2Xa
4kYKtfn2oxRWuARxb5SSH22jOv/P5LO8j0JuNM5ehTKFGYpYv++qKrPjoOrAkjNe
HEjn0Cjq3gZwzVLL7+brUWyE928v5NOyGb0mzHgBKW5cmB44VMHnU2TFduGC6kVG
RcAOJLk/sVF0tUyEKrGieNzmxPq1Lllne+GftjXMZJPGi4lyVehePoZHAD/DilPF
/qjlFKhI5b7+AqL1jlRdiXq4dtcnxrw7suIvCzYFwDXuttt6Y8o0SJovi/xOca/q
JH3gjg42XkEnaC8AZntMJiPLficQ5kC6dcQhR6/ZsJHgjhcVZHIi8ZYnO3jB+GgN
q7l3Z3wgmj2Kl0osKs9Y6Xt2lNuoYJqre1cK1Vgp+PBYr3A6w2LvfS0rHJmkv+wL
r6YbLdOAeB4X/6UNEORvRPdA7LzB0FqFVFDNwfVpXEUedPeNKh3gknwUdJs0Pe8O
UePIm2OeiXmwnBI4CmArRVzisHl4T6OVzPOykw6o5lshmnA5hfPQPpNHMvarxXwQ
dmNfKBjne/oP4puyfLZBjs6ouz+sYwuqmcxae79oGxvPmEtKeiAV2H7NQnwcuVmm
XPaMxp/ivdz4Wj8s8wkvZj+5Rhb9NZVOi8YIvbnI2iVyKagza5xCif8PiBh4Rwl1
Tr6sNshd4K04fKFSNKpv2c0QOPTMEXBCWFg3mM99xw0kezlMLrtDRhhn6DjDpKo4
IzYnR2LkOnaUWHjV0xdgOsra+zT8f3eZFC5SL1Y6p1XzzwtnNIoXtH4FPwmBCYKN
X3syj56l1AH66VEkdp6XRzVyqRNKA8haPFI8DC0/bZRGgtB3KQWO7JhXVGyooUgI
CvY9ABYczZlYqzNBnm9trb4yywoYvJFIWlJ7noiSwmkgT4b0B61hcay4W1fb+dtN
zoRbNZs3Tdv3xMvdx9tzorMKaTJQq5N3ZVdDixWl1bebUA2/dAIX1c+SbAAkbhYb
YKgR3ZySpeGixjvlqumNelsObF/217KWodERm3lv87D9JkwbsBpo/1vj3uOzm6TP
+OI1lX9SEWjsIcyENBNOjSS1CIKoJEbbaCBrplbva4DhfVAi1K9fiTQ6o67pv3l5
sg6ytksb6Isz9l+Nva6Cw76VvJMxyzq8Rsa9tZ0nsefe9rVJ8nDUtDnArVrJoDSM
/Dg3g5WiMFU0/n1vCdqBKp9NqwWq38rYdKZhH6Exvgyso6JE4qHhNPC4biSYXAyL
vcsQNFHP4Z+pDtaqPtcrvwWan2yJndR35F3S8cdg76Kk6Im0LEpYK/uaVbfUMxX2
DCb5etC9S92m8x78ZAelXH7ct0DKToQJHkaoyiacKfC4/z8AhpczAYxeZLipZL5V
Na/AXDFNkfkq+uYGCnaaAIeokRstxwMWsfByfzngvOxs41ePkOfLl20zcOHUmie9
jMo4+PHSbaDZyrZZButl0PgcyF0OT/3S7GqwqbGXd4N+x49zhKbaULfgQM8mvHXl
YfDG4X2GtGhLviExtSBjxEI+P2aW7pKOwLOHVLPjCZjy0OhYIVwkyyuJN50usMZP
WRvKQm+4rI9QX5+tqzezFruMYHc79KAoljvOAm8E2qvRNHkLQpuzBCRsN2ZDtLfD
tw/3yzoRZIi9qHfC6N+rY/I0ZYcNFrnSsievvVIUK3dbQAIWLjZztV8hA/EHqIeR
9BX91sVYrDE4Rvsm9f7Waede8eyv/L4wqDUKOZtIxtjZOQwgBUCtMUe+oLrFhKcB
vNn33Dh9H4wMJStAY1dIHtR57H1Pu/KRNbheH79ClN9mBGUtGTEU3fXjXo2Kw0L7
Hw5AX3vkXWOMY4aAof2XAhlbftiu3U6GSvHmpwl4p3uA0s+WrkxZ+keVPz47sl3x
tAttMm/FW0igkpSG+fwA4QVunTr0gOm6djm2687scDupTrU0BI6m4ERbjNuS2w0s
APGb+TLBwpgbQG6esB8Q8w2vnQ6xPxgH9iSfJLBNOZ8d5uFJV8W1toqHJDYWtN91
wWq6+6gzrcQoxYzaqRkBr99pE+xVFmBoi+sdWJ4aH9SjGe1CPGXKJvEw4xEnJawn
DTsygAxopW9aAeOLEqwBkzSWtYEmzZxlNMZ814hy23WdOZKx/mnEpXT5u4e2Q8vF
geOu0crY7s2nE6zEjJ/3g7m+iuK6Gd3n7To4l4W+tHmGliPut+1ahDBJvl3o5wnT
gy0Pq8RCC9x/TxJUovGnNcQETcj6rnf8Oqe/tJpD5xuWSwxAqifjRwnWP0Y2YOpl
BjucreZaOARN4oMNb3LxMriS7bzWxi7HcmbshMKl4Hj7ku40Zi16suLH0WWgordu
yH77VSxGwgh/9/ohrJQUxgyreQHsu1jiOXtBaZD23Sgy/xQhoiMq23li70K2gz49
ZRfMBMuHJokigUdIOawnqid85FBaHMFr8l9Vhar/78Ofdy3Pishfeh8gSAd5H2qV
nkNX7XFb7YzkM09G8VM992f7pv3IeTKBUlbI7fEV8TztSp7OWwpUIMHXzsYxCDMT
JyNgLIukBlaZdcANwp5+yDdmN9xUjbB5M3Jkol9uZLFVnQuSGUjz2QcIknmloGmb
XeE1Kj2wa0fy5NNRSRvppmeXi5+hviv0NFR2BoKC4AVIS9Oh0/SukJ/9JZ5LeE9G
uQ5sKPX+bmUlW5htNt6DyZWLKKMLEtuUxA0FmLzyQOsktI0huM2k+V3Kov6VINCV
hqLvToF6RPRIHmhF5+YsVqQvHThyAEQhDnkbGH7FkluM7DoGBJypBc0J2qAdoMDQ
wE+O37EOD8SNBJ07lrgRkYSGiZ667dZ78WPdzdfhgHAJcbfwGK41yFcRvwfcn/oi
iQexM5YWuoeEGOPc3mrziKhZHDjBx3YHKHXaw12MkxgiccT27vvA9BRU/LEFOLot
2MHlajq3o3Cj9Q47MymKNQL5p1seN0xrFUwVTvv21xChNGX1UR9fPycKXBOJNbGd
50rFqv6NphXozaMr5xzEPr/4FPen18SO5tlFniMuo+mpwgNfHLjCJcpeuFMRlNup
kNp24cOxbcokRJnOC1gc4WP1XrbBVFSrZ3RwE42SD7UNygNSGxlK3a1tk4Vnu4N8
H/9Rvacqi5eniqTEdTiKVM4xhHW9CFz+tYeWBoaRsOy+xnZjiGzDoatB6lNqe93U
RGQWNDmeaeVmLZ5Q1z06HM7n4ApirXFnVKPdw591Tq9jTlVV9hG6603CHy8IyAaV
GoLQ6ZBYaVabW0Ve6OEA8r92xLD/RE9MXbcjiAVA3mDhyB/lvnVTejxve8SKIGti
e4GZR9PCv3zNBqek+AP2lKw1X5GGtO6qYAiAtneSmuGMcqjGfItEmJ0zHPpzzXPJ
RxxybjixdY+4ep3/qoo8Psk5ejRorsirTk7JtW93NWb8thAKUkso3N/i6RsMB0j2
WSw6u+WSFYIbE9v42KgcwUFct2tAwPB23fYVF63I6WRv0yKIMY2Y5tlBHJsyXrFK
L8DdW3aJ1OzmvRrE8GO5jCYmZJo0vuYMuYZTzRR89dIRAqFPWghwOcjZp8LJuGN9
LgK740atUkR8t/uli8gGf2K0kce3cMgd8QIhuD4GSU53GcYCXOZeMhCEAcjopC16
bqGdWeNZJoMBQEdtYQlinXX/u73psfjr/rXS036ZKnfwMJ3TXg5e7ZhnyczNdrLK
1nEPylaiAjacKc0GbBE8NCF/9AQqeFSxszbB9deebsVbqIVlRMEXqPMDpwvcFtIc
vVxC5O8vxMmZxM3W1FnkwXGdiLiStflFNB24VXdaYnljsOC9dXCq0O/gROP3KHtr
FwnBorcC+wDNWDPK3N0TUkO46+fT5cnpiAWYy/JsikD1+Y8dlQmiUp7xxULGBuaa
xQa8Io3XpMggaFnWX2VJ1ogZ7Qa0QVjDVHeaEyAqh948BdAaqvtnQsC9epglDnS8
JqlIHqEH0/f9KSUdbUKQNLc83ef2UzxC83UD7UU3BWTxeB0+a4r7sp48KrnY5XrT
wD0XuBRrDr+lyf4JSMCpL+W8MlU6WTJC8IRHdfilEPC2LU0kEI93ufMY6KE/lJ8b
1ynGivwurZKZXWnGTb+AiLqJawzEawRc6FfIb4cB2w9qhMcSqEh2Vx46/dgVfzNh
QM3vVqsY0kFpDhlddcuMU665cdTfX1a93BK1uwNVTgA6VC8u3NzVnzt5E90p/Cmc
oabAMJ6OaXOApAY3Ezm2TIv+hbir//OMYnWAv9AkOCtrfhVd8PNirQflsHKuZgcI
8+ZhkIy8RTIe9rC/ZB1BbEKSy+fVY7BTSbG1GE2beAZ4tDWUiQ4PYLorAmn3ygo1
XODdKjJq8cw0xVqnTagPrapG0KgRdak2w8aoukBq5Mxy+yvXAOJpJsqVyv81npno
KSzENEXHvQTbk8eOvYU2LhVPq7sIugureUr6CpSetsdpJmSBRyo2ruNDEg/MhwKB
xdxMgAyXlV+LR+mPfYWJRl2aVUlmFhCjMhKbKGsaWhrCFTqhhm371E7Y/KTXWWW0
VjmPcVk4xrcYXNr1W/MGZ6rkSzoNpskisybE8ANmpv0uVID8rtFQVd5YbAtmMVzL
ctq6sj5gYrLekke7r1ov3rRUdeCyFN4getSOhRqpYzfbodG9sa9ZCiP0SSjXIGVh
IzrOk0fJ8tb+xMUU9YQEGsgC2V4Q3veWaMsW6Qjfjiuo1Ye0RS84YyuyfaqcCusX
uj9i5MS99yD4BuM2Wioq8K7mpqt+ls1ra6RvdMUysd0F165EVMhU9uC4qz7ri7mb
PGaRRVBCNvZSKu3bMu3aP9/X2ZFdOXesF7tz+sQ9eHE2AF5Yd1DeBM11sys1mx2X
+DVFAu0WP7vgSgMcEK+iE5VqZUpEkjt1iB895nCWNv4+puByDHTwLCLrJrA/xQ4d
tx4Cw6nXhKc4fbhgVm/z+oSLgZJrMm0cXL6FK14929tREzbigfRvv/KaXB2iuLYb
7HFwVzNGBQQrrGhW6TAni9sig4K0pRk5n9rcDRaOPVd4v/BtKQjYKrXGIuFejmh6
JL/FuNMkI9O6yGSyBBjb24NEMUKPMgTGbj1vWlDMhzy3H7cxw2WL0u352koR6n/f
+qO54OTlFbOcDgtN93BEZy7BmBvLVP4zvIRWRwKk+2BsM1nh5oAktIPqQJNJwjz6
M8AwMoqPmEDrWOLv/uNZOKU2158NcBrNQQ1FwetGUzeLFEfZN8d+YvSm+7PZ0Q/L
T8uvWyL2hghraLe0hAVJb5G1MBmhdz21hVwRJFtiwI5H1v1oR1mwfyUrILdW1JI1
8HLHCWrcygzFjI0LSa/ajS2M422RCxLu6HoBsU4Maw5p4E/1Uc6A7sEgrSFDn0TK
JNUoPX8EmaO9bKIGBsR4nGP3rK1aD6umrVR2w+ZMTpP7+hGIFd2LaBm8ltCoS+UD
dufLNygQxZQcL4yDStRv3WWAGfwzd3j8d93Z9RP34f/c0Bbjo2mlnuslxovd1npx
PR9q1LOadBExdWcOkFdIgcVHDUHDUurLcDs1n5bdADK00rWkhFzo1DHs0JA/VsGT
cbUCIy38p8QaIDdTFSMle9AVB22tivPcgekAbbOZ23yqpGdM0ovORe3bBdUd/GKd
8uq8RA6OdvNcMPJYWpar1ZkOBCzgxbIz2qUgNkIAy78lzGVp+H7FNnbnMs92odLr
ueAnafYxebB/PiuSVmITzG1KUg3WY+tq0Ik8YrlvtJ5GgM6180tEHgJ4Y9jd1MK9
+/BHQBCctZTR8mE8SphOnl5OrGRn+PoVPMwhJuPAjCj6awIYndvcTC0oIwQSgldt
UvZyMu7haBryZZeUP3z4GzdJ+tKvqAYaBlXr3rAxRum+MeON7mIV0nhDwoYisgKt
uAqwpkOB+POY+NW3KRsGXjAlObFO3S/RdcrR//nqM6s75MkPRzEhyGTsrMHhZZwS
txHdU+24IxyhsRbTikL5AO8ipqNwkTdCVrSDDulc38O/h0H44gKKquHD5rsEb8AS
85E44fd0qAi7gx/RlGq0qPLzNaWRC8Ym90Z/9AYzSuUezoSBMsJS5VSl9zFyFyF8
ypTBBNl36Yi1PYEp/B0DakEQIG38NmEQ8Ld5s0twHUL4BmMe3uc9UZKmgEJUXGoY
ko2p1cWOj8Sp4IVjr49oNG2RCZ9LxlLT77jhGi4H7aRsmFEULT097d2dH59qLtBM
uylsviVXOcqw8EkdonbKQ76gie14o0L6M1hX32O2qHvRQDABa3ijNLOgLyXd1L3j
ijW/eO5lhO1jTClpF/7Xu/t+9XAmfCZctcadLIpJtjJkIbeZaz46/Yo4WSStnVL8
t2E1hSx1WFL8Rva/6WnBM0QmlVNTbHVWP2LD/7ye/3pYCXBCFWWGVlBT8aMmuFfJ
THXogn/PuvsNuO2O83mUuW1SrGo1IbKp47m4RWGvQmr2P1e31aQH0TKgusAss/+h
atJr5vuw+jfDsvbqCy1yvC4qZE59zp6bvjJ1qFsW6cKlhlBeN+oOsQCGFYyBIoaB
w226jbplzBjQ5q6Es5n8zHnBUMU5+cNUlr4AAlyQLXtaiFNuCcN19d9xBjl33Iga
7D0v2D1JBV8myAHoOQU+vL45w8MFv8UV512MJiyvdyasnYennxbLO9q87RUSG5nF
jRXykbqIxfjd+cDDzvd8uY6Iq+p2qLx/2XjmD8V8XgkA7m1Af9RonZBfZlCscdTJ
xrn4wMdTUykEhiumEXgV5G5b/6p1uEaeVjwHF5mC6iHgeGuY6EVzO/Nak+W7u6M1
k4WAqGCa1iKVRzj0r87TILIhnfnYsxVGhMP7R6jeJxa/v/+vLzvTlfkb5ceKnFUB
G/EFkla299ZD+SNJtNpwQv9j7/HNtRZRx/o/+uLh3TFI+fZJWrBMqRGCREoDPxKC
nXAbjt9CCyPQcsNbGXcclfyY2eoundYRBgvg5AQlbUvt4Bz1y9wTNAeprJPfF93p
3LGsyVP9fwfODv2c5aEUaOZp1eH2aOeZouT/5S+BrLV29g00paPCHKePByOaPG8H
KEc3bneOOUPVCMSKa+pgWr1qcNZWrcD82axVqaDHofKBvCSkwx5tlb4whimTHbZx
AwZSN9oSefFHb1npcBLVlFMCL/34uOhfwYwlH61WPPpvMqWjzw3afUKUit5e1/rD
WGLIztYDZbyLoDw665yh9KpyB00qVLuFIfFxIha5rlqAZXPQC0F/RNUYU7/WJ3h+
mfRHVvCkwosghKr1+vqXhcosyFpsAOEtqPvYaU/YBAChvIck3XpRBXIhbOUC4k9T
XXJgwPU/ZvA9mCqWXPQ91T7ekG1SxmduqCHHIqtqj5vdtDoBYWTcFyZphcArUh/N
OEYTjB2OY2GpubQhe7udx3Ggx94pDXXohYB412H28w1q0hFpySXXDcdpkmE2kgqH
0bgmUYGaLhqb5zYGNbIq4ftCWpIdzRgdyrSLt+bIOu/4BMZGfQ9xKv+k/fTcKXTf
vo/U7eE3BZfjQRHFD7vJ/7g/KWnxq+osBT7NpPEU/arRmYsalKOmrnvP7RIRiOi3
qdA9ODlIjaZ7g8ScRbe7+Fsq7QA45pxo428yExoA055X9yiHiCur+jcVmEhPrmtY
di8/HSW9qC1+4VO0PO48p/P7X5DCa/3VijlHJhDgd3pxW7tfsM0zT414ec/daR7N
J+IbcRQqgWaLM8HaL3MR+dEY7XLzkWuEj3QJg7BgftmuHsczgDPw8IPpMttwMQGL
E+GtsUMNuJ0qCbkeBOh7He/GTclM9JkYx0UlYMmmrn383mo5hal5I8fpaJso+FpU
gTDj0qM3WKdnu1yis7KMuv/ucimAZCbdtlQaK0IMgbczx8+2RyznyQIDJy32aLqJ
ozPrpT2BllC+iE8j+pAvYkHXYzX6M/94RfWMoGc/95GvXhclV/UAZKXAG2DqVXkb
hFTr83NRaP06D4UtL42wwTw7qAG/hEl3U05lhImdIaLMPxcCa+0CP+YvlRC+NHl7
pPdRJVHM8S2xEwfBcY0DX7+T1VI0SU04gUP5nscSCCx0HgDuHuulCq66SCn4VYl4
sY+bNieNO5ld/S4ubKH7gwVCjsNhh58Y2n2yy37We5CoKowhbVa+tXKlu3CEZ5q6
O5JaZh5bZq1OlHX6h0Y6E3fOQoZPDumntX2bbkhSe0JeQRWfu74d/T0L9es3p72M
z8Dfxchn8CWd/59qrdmD9ANGS7W52tAINvuURli2Svx1mSo2c/7A6taqA3Dni2rZ
ztEpJmVtGN4AHcEpyqPBqkzz1rlPzigq8yMF0F9A/82aomv0zUOm3m3gyeUhiPF9
66EvWygW5WAs3lioX2tcrcQv+Rcd8MyYBvesiG5FG38El11Zc0dWDP2JhgGBSFEm
C8fS9bBlKlZyYhI+NogtfGjEJoNeP4FtchEWvm1QxclzgWV+q4yn2ysPQtt6TVV9
chiQMIaNcm1OYznzrEMftK/saGRZqFJQw3Pb2cKmxqOcAy6KRtMClJU9TaGc1ZFM
m0XMrlBYe52rkp3fI75YbxAEoQ1cgpIMyZBbvAE8x2n2AeuM+BnMoW+HhY0/40m2
si/r2Vinga+EHnCZ4xea+xR3Nxb8geonTdN9ZVwSpyBrb+mVH5/iHx1Ht+FaOSx/
IhPVawTWHpzt44TKZE1iZ14PYLS24mF+kvKuVjilUA+Hbf7CMkr5B0X+XKPWLkeL
BNyDFEugFWkXjdyJpOD4c4nRbE2R0fLz67XVHrXYGWVZX+uiYPNClcR4t5447tO2
hmiZ2mOFa+GbAbCjGKP3TvxUXNK7pxcVAocKgualXupb6PCz2/1F2JNvealoFl5P
cxgACsbM1TE0h+V8ZzGbRQsKFSccPezkD86BnBQ0fak9V5c/Z6LCC9v5u846yCnd
33oIyJJZoO7jYM6nxM+65SOmaEfvzOUTZw8CUDbwZiX5EBgT1e9URWhVzaTZOaJ0
PWF2CWzOjToIHdejegglP0A58MpplZE4eEn9VmtyjpLWLVAiw2O3joHS20+ZCv7J
EMrEVQLbFp+TjrIt7bIGf0bcsduNBS57MwO35o9XL6ozkXoPEkkk6aMVkP3EcwR/
Qt7nhIPubNg6F0gEYSoUBhz1lsrj6XeGAI8XPDeBesvzRxzlwVF+261UzMcMnjTU
DvuABckNF2PCJHQcudBCrZ4NmWYwYaZLpAZgtpTk7my5/XX5bFfqL03D4navuAzJ
Q3UcBdOwim/RYUrMO28RwIh7vmgp/4EkUYmTaOqnHiF+Vk6sUUdDQDs7pJw/DtU5
LAIv9RzpUhjcuvRAdLFXn2sgQsHC6KYkIOevtU2t5aF8gg10wlbChX6sdXFqvaPw
rJGVhwv2vqJRQ2o6xf6QaNkVYm2ZrePgH13uiIZGLfqS3+Z6Ax9P5yJxTatRJ9yu
sojgxh5iTwXG/IVfpIzSR+KgFTbTyw6Bw0akCZxz0fOGJEnDZ1Rq4GP7ZMuXGI3s
27Ha8GqRaCoVx+YW/dvgNNp0uG7JCaruQiLfuLZDtH/dwbxzEqjvrDLn+IB/PhF4
/rD8Dw1Vx3W+iRRxgFzFInrROr5zPdoI0KS77hfRWHgQ95fbBhXuldlhqBioU3HB
CNv98AdEYSfjXtW9MU4fryDNM6yCZTI/D9iAUcDmYCU6Tk9/H7pKi6aFkFkItbYy
mepDgNqZitGdqJJXx4LOkAh5o/4WDFh7OQ0+K/RH04C1JGUqnHy25wxWdmso7k3N
pfzUk51EkSJZ/LNtm5Aa3EHrPHS7sMlHm64qfA2aTVSZwBL85JSj1/VPzxjms64C
GpD7fwEQe3o6ELbdRBjxaSniIgZOxwMYMUz0rScf3dtnHg0b0mtvabpgQVbu6IJg
cNXM2KueUkBvyeDrcmrctF3uPjIuJqxKsbqQm2wIuIbSwCxClKoxR0OBkiN+niv8
938IXJ8+JtKSMyp+6m/O3WnMkfjYYOWw9tL2/+tfjAtU7mc6MX0toJPpnFpnb7le
/xGiyi+eUNXZSOzJ/vJkp1wAIijLQFbDkVRrHACmKv6xQL70sAe0fmlPl1qo4nBb
d0RijfdCDS8JjjZt5u8N/Ft25KVhhMGJ5LXaJ4ppCsZrMzrB1NVPnbZLN0yko+gw
9L8tcWhHTmgmmE/Fplkbeb0Vttc9OD9eAhoOfWAB0B3s1WJMRoKzIju3cbAy8tcA
PLBk2h8kFGWAkTNQqkrT0xD253/Qw8Bg6guGXmvfD64tM/Nmdr8enqjmLZCoQvuT
FqxWBrdvhd7EejBjxpfszGWt6r2+jSVMTDzLC4/wO7X/NhWz2vOq9cnfC5i1Asvt
aCCCju9oC6wimlG1L5r3nn4JMR7mttaWOJyMiZmRuOXMXVfQalrOoH+1nbn7pag8
ef218TYrEQj9/GJ2h2rHGtb83YFva3qFUgxwf7OKiRKzC+gpjWjOqprgjr9Ib5yC
HcqDiPF5yOyZkvsEpeok+th3wE3Gd6qEi9CEME3ysBuEzz7kfmFk00PYtaDreEK7
oq76zAqAClOSkM+KvkPBz0wDp1erTXMaom0W6D8ZIQXTEdahoWAy+0cLZJ36N7c0
Feld4mWnuGUhqBIrLVOIXczGwXHPsWvlZSuHSDLqlA3nVkoa5P3sl90KPVOzXAno
Ds/zJeg/OywzM93vSCPTBJWsXmbq5xOoVdu6U6gvsXhbx1gZS4AgvEe1dFwUGIJD
/I7zROgqNtWJhyaRmbgptGhl9ZNSdxpug1m3BVRBg3VTXYAYF3wrW2lWtCxMiNC2
0iGiO1RikgJA+7+ehWhWN/wGhcHuz+pueUPaKzF6YAxY5KztHWp8+MYH4puixjFV
GZAOG8am2/EafjiK6bbjxu6LX4sbz8KulJ6/8XAl5PwXDyXgsKp15Mmq4UyhQSPb
vshc6gsS/SZmdiLaKJxGJvWWQ+ub3Mc3g90hWbhBmrm951gHZrhPe9hLsklYJKPl
OjpBt2zZMAwiJn5FQh+2/BxYxjHNDG9CEmQ4AxQxXk3n+xD0eAVypgvtJQ34+kFs
rp02NfIZ4ggUsej4YlXm0mw8tCWrsii+fwD6Ew2cZHIsPOdbXvi2L699t7jfISBV
PYzny1DOPzvDLNqs9xya9pJCWyiBm/lwbASAk6VbSjoTpZ1MD7YGJDfto1u6ekW9
97ipj7SDRIs0rSwzvngcWvNJMck7GOVsKKpvsOStIIWtgAZsPLI3Aua4XacOnTNV
EVydQq2gdAqVNYkG45TLLZQ5XgPA8Fde+Qc95OQFdP5WmgqxWR5DkRFJwPsUwnva
5XRX57bG4uMgQz5otk24kRRwWmhSsX64r/1OtGCT/WmSmtm0A9MdkHWdylkQqy43
LDxAudrvGdLd8dPp07w0caAQ2unUH/gem/DEDDyxHnhB+SGj5MUHv6/qPkg1WW10
BlVBa0aI7B96JEwGgKGX0WLmOChhN0dLuT3ZtdE0z85QghdEuV76AdURGWK37XnA
DOaU1ZPOT/UPIJgaT2F5AqYJOvX3SouisGCfnOwC0aNMcKKF0Ix7lAf4I/kCmvuc
KtxEttKu7zLYd4LoVj8vOHeJzTzSfqkdVT293P2mP+gOJwftgXvZzDhJeM+/366w
eG/Vly42LPoSuMetPRTYMTlACbZ1k3lz/TRyFYLyak9zLefMnpTXsPSmgJrddEAQ
G3goEKXhW4/862fSzmDD6Fdb8DAO9z2xdt6pVLEhKNR84uAngen/NPmpyQar4mGE
s7RKGD+MaT1T/6nHVCL5sM620fgIwUM2IJKohn6bqxVrHBUkuFI2K0hTVr3K6Jvl
OM7Xin3WpmQME1VHorVURYJNgjTQmim2C766YxZMt6QWIenHuv8ES6hJJ+dpEs7x
oF+Xu9f/BXl61hLKlLOGgj+7kKeaHtEbHs0lQbVIRSu7WMFEXiHFJBh+AylInN/d
NljpOx28/4V8DLKqsdGgO7JDYCCfvdFBo9iw4eXi7IwQZpATtUlL9MA8cZ2WRxmc
+13K0ad0ud4KfO2W8QEYyKrULi39jnrEyXpk9Liee8Ft85Gpd6Z5wUWY8EoEP1TE
1TgsmprIemiVZCGjihepDTRNUl20MIxsSTIfo17IXAiPUl7OrvXTxg7oEtGji32I
inWtrW9Cw92FuAg7967Hm5VsT2np9of2y+E5xkV0As2Vh0mGaXZOmFzkx55+QdJD
b66ombRsIZA0lCk2Jy+M+oFUpusq6dLQYRXfMoseg4ImjL9Mlpbf5o91ZbhdqmAg
Yky3c7LKppS4EMZJ1WUAF7cdyCQr6+tc7cqLIzixRrNGsRR6d9x3TDOVUX6FXfV1
KvArWvFMr7wPiWfKNPHNUomtcVMYyFfWa4Gg/k7JNi0WJloG5fEt7ESZ3DFcs6Em
fi5uoO7BnuguKiu0s6K0bJPWOJPDJKmB4H1LIv9RpDP6W98/3iIPL15rFRwOTgjN
j+wrdXcEODKkHMyhmE61Hz4bquioZVwS5GUeGzQlWq5xiPC45HCWMiKCHi8nKPOW
4YIFGRHL/FDN2FHYOw9BSi+qotcLd8JmRMVAKK1GA+O/VmnoqhgvHY5U5dkqtl+r
quDNvZPj1kbUiUs6MbNDP5yLXb/bH3IG6CsurrySZa1qSyfuX5m2g7cDP9i7tMyk
ouOOQq+bOH/63cQQxtfG1TLxmHZmgLCUeUXK4AitZenPU3FbO1vxuxhOL2MLL8Fy
ZTh8NyTCa2uLbLmx8woAQQOCY4d43sU/Ypq51io4MthSnpJR1WPFGoeNrQj8/gEw
lUZlPtKdHrjmJfjKuqLdeDKZxIbeeZs90+6tqphQnAgy+yTYmNikkPhZlwErT91Z
LcU1xFNj+JnA4sKv9VomY54IRui8J7u6ub4cK6biXyNU1Zukutsn2YGekcuQKQnQ
/Sn6Z4+eYtVupseYzPz9NWiV5uocUV2mY3QQ/9S0GDSaI/BgNpH9GQBHsrd/O4NQ
MLke+4+YeOyr3zBpHk3gqnO8314fD/GINvmDx1mGlE/PjvPZ4i8lm/PkniTwgT5J
f/O4x6fxoKzNc7VvLVfbIK2CpUVUuJWL0SBPVysX8SxGFHTe/luiNuXv4GANnvry
lSGUEsyZzgdV4M6/rmbcA53EXBdutib+qeMcc55KdhBVyapWY+ENyA4+n5Eh+fFn
SeIgOJ3wQOnUFWmzaTQGVkA4JsiyeyqZhNsAicsFE+D2L4fS//oKIc07oSlN3oSQ
Po4Ub5Z0oZwqNUp2zdC9Efyo1NveenQW2z68BUsfOEXlzVzYNVC880CQFPw5/UA3
gkhN0cRXoiDUoUVXts08xrTjF0OKoPP9OLYi81cMkoRpb/wCn0vdOZ4LF8cBIHfW
WIVF6VRykK7BjwBY0Cxz9Of+fDJV4irIWF5ynwOckv1YedPjvgNrgfdnLVcF6jZA
YPHD4idAl5xmTsWxiDoO06q6PhFLMtozsBfcjTrvZuUjdVUq2eZxR0+t2XITUiPX
fiqoGZqJWmvJ2t1Cn/uom/lD/vLe4j1HUtkdaQWVXLqV6HAERbrPdbEbPe/wg3KX
UJsQi7wCHN/uYDy/HlOTseef+KxQy7EnhdaHGmS52Aao+y0LBmzAVoaizys/heBN
ERDM13qhrbXAtyeKUkYhCPjpmCBjpayHW3fyiFx7JGnZMhUDVvUXU0S8RZLavWQq
YXe856zSEllCUzRKqVEDbbOmLjhqwrdyaGcdr7/XX9tvwRogzIq2jxZ5Ts2fuoMT
dSmBU/eNIHdYqezUDgVrSUSxfXtekOKjoXpf59RcUAiaJw2eNvI5KLqh3tqSqcj8
LDSOs9NYaCZNxoqd/IbPyMTloAx/5+DLZLoaTAdYnLnd7B2abJlbZqH14JU8gHZr
orZdTq075ZfC2AY7Y6oRetCQIWUsq7i2Q3obIf3DMlC8eNcUS0OBsLB087vxN/bB
dzNquQD3NuuMq0/kWZ7iVrVTsy2ncojwacyfNtuCkjyg2lgIAAXIW0aYt8jpRNUU
dEKTglCcqVxGRT2WpTQCkTvNGOXhM/kltK0026Gu3plBzJ5qVBYYjbKk8omg0WmV
WNcYHZx6Cpbvv6aXoSYKA3ZOZ5dikD3ymelZ/CLH8Alc8oGDPbz9ayRwNym1+IeP
YCWAn824/YqoejbQL7zoBWrxfSJRdNTXjipeS4GtZrqWKqD+18cRhLxrYUtr7J8H
BHjQQCIKEwLCP8FLdXi9hYUpNnzqeGM7Ks4KkmUl3fVHfp77rdSCkDSXZCwiDku1
YiG7jT8Abh7m1gVMKbzTDb0MpIfmNY/xU6h+KUIUFwjlOP89nXgKvWUnHhrrwJrp
AfHIjymgUSrwKdwog+JeiTlm9Fo6ngJR64KQSY+PFkcWY/wIZ2i91iRYlb7jDD4n
13Xk6CC8mB7wRXkCC841C5k36E9H0LE/3ufY1ODO8CT9B9OIsob7lJ9s8Y2rzrrX
DAiTOxbBYpkb7VlWUKxSqUG5C/i+DsPqmlVWrX1W5Zr1W+1JtmbSdoV4nnU+adZq
3rl0AEKbfJzYsGyUZ0GtXM31OTnXc5DNOB/fmY55iabhJr6M02Dr6Yv8rcmE2Ovl
MeLbxzQXyzSx2XcBqSA5PPFGAwHfoDR3wFgKnNSmEaFt3S1WijBWiYrd5ISucTha
hK+QTj8W5Blu8QSx7Ah+86SBrfnGAAIGiKcWVacvOyI3VIWbZiF1mOs1K+rr2PzQ
r/JTpaJ74T6kZ/AKgprDZugSXzqHxt6L+mOwrrATdnKzuSxi3qRgpkIpP8DlF11x
oBxj/+5p24Pz84h9BER//5l814SszLMXoNreGRwBbtX8mWMz91uuUDBvOw0RFM+f
vwjldBVHCOSr6GdudCo9a4dzSyLNI3ShS2cr/TcUVJzQHEzMDY7cb3zkDqcnW0dc
6Jiidz9KGlUBkgJtiDpTT/g0qT1zLGqCJnbkN1s52KyVpO3aYt2Ta92ZpNvjtJbz
E3sxqZlQP3Krzk3lXFmkMdkLvkcasklwlVvALFR10xx47G/KdyUuNs3J1jLhjKM0
fND8F8aTqaqohr7Cd776b41siZYqMR5coLoEJZb9tTdjJ6qVry4ZQyuV1q3IIHxt
Ka4SYTHVnsZhyoPqLfIzBLEl7vw3/qgO2L8MMyceyQhMCima1gV26kEnAQi8hE4M
Ujaos8x9P1npTTbT26GJitYnACvq10lb2aOjqTZTDe4iozfr2F5nHr2VIVc0ZbyF
FBZFPo2GVkJCU7FYrNvoVZDtdntT0wwgNY5ep8c9Y5vB7uGPHp2a6Kvb8bByHgMj
k8brvJqB68dyxDkQj5a+nFoO3CrDFEkY5JDsuIddltDxI/ztPii6eMFTcsIQjuqY
bKmUT7WC4dUc7UjlMjj0QcKGcZ5wjk81iQ6rJq/gu4rOfRkZ+3dHccffsebbo9oQ
/i/ea/RHZ6I2DF1NBX15aIOst1GFVrJxnjTMGdiQIZ80b6Sz6X3DdS4v9GjShZ+t
TTJW1YLLU+MUjsNhHlRt3xI13jTodA7R1aG1OML+/yVZwpenH1XUDMBWDhB5FoR5
0khKHBR3qgPlqNmB6fxBmGaoPC1SekhUWy8RXuhzEJ7sU3M7ivS8g9brR+TBSjWq
GSFdOSjtbQlGE+UkxPtPcY3ENigA58qEy7Ej484anLnN//tY8pn0YUgTzeeJeM0/
wW72TTivLco0lbFJt9HFk9UV8Pd/iEKPBI8Rh2qTQ5vQbfIW9ajeHTntTyuh+iVO
aRKTBmCIDSv/KOEGLJjgyfEphFeaC13bqKycsM5sKUosWEC35xD/JhvLmqcFdQUB
3SP7wHSC3mvhjEPLCHml8uebJGNxSwHudBsScFsgG03LAFUVviyI02iwWGIWqTlf
YT/l5WoDDyk+tC3XbTSuLEIrQ1g4vWJ4qdygV0f48Fj6mnIKR5ohvEUniQiHNwNH
T5rRur58LSzTVY8SEAlHtGOusOJXv2kw0+d8RZujyBWtWkQ8IlsNtklYZeWgenUd
B2ZZ02B2CuxoWblAphfmocPZWZkVyf3N7fwZLmdsiL2+rfTPpsp6i/FOzPxiNrzH
Xg6kfFtDgrjfp1Zn/UJJT6nx8hrZgb2r92v0pPLc3P8uuLjirrveb9mugbMEsdo7
PWdOVqzNjdkBItDMl7cN8pkIpc2ZvoPJBbbuRYl8Q+bXTawlDuK+F8Ox6CnIpmrZ
YIWyMWoKuYcRbU6Nfs6YDKEYNU6W3Vk1PqN2sqLy+fIQBhcP5uTdtmO26BZvteTu
lorw2+QaxhkX1eQcRqENi7kHdunOsjhroNjRgZXktUzCXJFrOUMg3wifu+mjRqS/
Yk3MbrjETJzDOn6NHtCjGAEB/G06d8N5uhUQLFqJ5quRDT8ijPbQDLUIDY5kYN71
/rGVm4RUzjbFYgQdwwCRmNKqoTacnosQliKdW+BdBsf/HOe7qScp6aeuwq1flMJo
yfYucWArduzwhkDSMcuHERxSGmPgH81DIlehTiET4LS7B3R5RHJIUo9oEf2KdgUH
mbp/eDCpBlRUn1KKuIJECDc89FZ6WSYkQcowjD4RX0yBHzSs3NFxx4PTHeRkL+/h
KUQUrJ8Kentk8rQGTBYX/L45KH/2PwS6/9pW3gvbadDrKfgkJROQV5c5z+n3vSZP
6iSk82gKGcvdIl4PBuZ51Z8ljJ7veVUfUQAG6+OXOU+/DUBfHAU6+t0zv2DqHOws
s5RiUePG91tu+rdO3917A3OQLOvONxT82p1HBJMKOUaao+RRZP0B5FnGJmLNoVjN
MQqaqcabcOlPCcaM4tnncPeuTrgThLk4nZSoRLH0VYYWzUX7Sd/MxIs2PKD9fcsg
4Q9WEgwMHMyBC1TQdGrvuA0heeJjIusAyF4CIkbXFfdPSNhvaZkvIBWP0Oa8aB4g
AsB/lslzXdVlrojMR7xSEz4RroQES68KF3CMUWbxoXD0/BRkeg/tCTxsVIjZ7S+q
nm8lqDv6JsavvNoFYN2wLI7a3tCvB26boioUGrovNy0Hu60aKyVb7BKeHxqhRCfd
dx6qirOBQz1+ZkeAaP4ogS6nYqsJTDzpSubpaZG/QRLeNwpW8Z/wH1S1qxREWKOP
LSI8dTRQf5xhrXlts0yy7oUo5C7JGgEqwayu+YqrbUSrgcAsnIwRnmW/mJAoQoqm
uY3d+QMx1KWnFxrx36l5aDzuHg+yM+clfvgb9sJsssBVHVbDsyrgf5h77jI3Dgjb
vINAUHLMzLTjkO1skTb1a8IojFdIp3Jfu9SQMAxHFjP62zYsAfKOY1jn4cjK1DVR
3hhxrSiBWcKkhHobo7Pi2mP3eO1nBcIsY467XryMjpmDZiPCnTEZVZSTfjJ29XNk
DjB6fGgfLX6RPRJGhfMVEVU+jXtLWPTVq1+7vKU0/Y9ihQfQFofYjXxmu7oDo9H1
QGZSuZoQvFtEv8bt3iNQZXZwtoyOUk/Ky2I73RGnUqkI9s1ag/NuzALJzNkD8L/j
/zM5kW4tid8l9agRP5Jr1QmOqV6V3R+Z4CrUp/9X68qnVsYNoPNoWIm4qTMc/At7
GY0VnRNfybXH2WmZ2T0ZTXLW9RX2wjEE6028eqTZHgaR55UqaL43Pqdl9zO/TPsB
61NAJpY/kjImEZ8vFZoNtGn5T18yLITzjLkGl1DkZ9P5oi9O5sGBi1/3+WUIb923
DOFhZVnmzhHAXWtkgqF0RJ+R9Ca5bDnj75+m6O+xd6+83AWz+yc4xU3xxycV2/Ae
s/T09G53S2uyKhKfGx5DKGzvoJsxOCebSJ+A6C/8vCBexpAWNzPTIVluVvYZw1gZ
GhtOj+4xtQQ8WjzFwQBs098upc5s4i6bXlsqopX4t3D8SDzg0moWVPkTQzFfi3QH
OaChX/8ceoav1u0a2fyAIrTpfbLjiK/U6UGr2S78qyiOPJOMRJHiJ8O/zFoHfkKq
uQ4eeT/Xg32z7DDDcduicMAoK0hPWuekP3ujXdR6NvuDWfF47FDEMX5cHIcxKLXu
EadJeRM2DHBPfVNK+/Ov2YhU4kffSILaMh/6M2cw1dEgHSO1iI1pQd8yH0ht/msD
W/wMI5rjZKELtOo6pbLR//p2gCRwlrbeOn7tsDra4BbjXVGKeZ3Pcnwy/vl1nAkz
j+IuPrqNil7ViPbEjERt9YvS+YCgiz93G550suRqOAh1lESzFcpyd3pfy3PYvHV3
Fh8hL2uEDKgkL1/uMWIGM/Y1AvDrR8kXvA7bMM9f4/aWoogBU9M5HBnnuIPu/UYw
nF9pYKD62M0cpyQU9AJkwkhXBhGT6mplusOjmpfUKcKf05ZdP8sHBiIVKOsu2+bu
/CQHOhdvL9JZ7DQs0z3XVSP2irZ09jfuup9Lv2SGmhhmRlou/EucGzezU3VDuu3R
AVG3dRyucA870NVHB4hwunccRoCtpYRGWP8tB0lSL7ZV8Bb9C26Z2wlmilEvP/J1
hBEa6pvCyLPyAWRcwECaU674WCw1lt5mUb5CTxGDug/wBn9xgR9xlKNa88cX78iG
9F6uc5mYO8bywPZDmzfJaJN0cS2sR8adqnEEJ5P8jihTtaQTnZq2F9MTJ6/fgRNy
HduYLSJFrgWli5bpb7mihCX9OayOpvcLqFKONCBUSjTS1iTunKEUKbERA9kPkFe9
PxG1lxk+OL0aMUapbHpypdvWxxKaIO8fn2ICA8JIDX0aYn91eQRnD8EH5/AV2bom
EOYSjdHiu7nYOd2N2IdapGybTraMhQlO75J6j2C/8UpPyjRFzayqmaoxKdzCeNdF
PQKwpahdpyaYDv67KSrg9HMyRiGe1Kc11nHCIEI27r0iD+myx/xwZVLV3ja6+W4j
GNEA9puYZ9/XnFj6qSKnHMtSBZqWSQzLw5rJInymfqFp33rkimr/P9ZmF+DmEM+/
1RrYk1pLozLlMwD/zzNp9PnndOFQCQBU72+im/JfHt3muQV4I8qKBFXvhO5BW1qC
p5zXhrrO5fteu/BRkFHOlKT6D8X6wlS7ZVrTflJxotRVdAysmh+cLd9D6h0N2ZG7
QvQ7M/qqL4tOq6CLy29iIak9Tqr37fGVXi2phdH6KA9V1hcJh7HvaLdef8t0eeQx
tmJWAhO+Ged1n3hbIRFYE8W/Ueqxx0k+xtpxJi1jTHnr4QtzRVMG8via7IStMna3
Kae+T/crLthyTTVC/SaWjXDzIkPnTE9E1ZydiTRiYuzcPPKj5E8fp07dRNS7Qscg
m7srbNJnLnadm/SchHU018AmAdeG0gyZBWdJ2ho05WQlM41M+1GN7XOG+OWX/Ftg
5JoE8fdMnDNcL/dQoi/uxQiulBUxQlDcHmi3OVkL2nuIR6GtP7jp+XDlhzjg+AO7
6J35rDylwMFC6CohT9mfnJp98DhMiI8fSt5Qe44dFYPxagaG4zzsjzJuGExsSslM
AGLKEaLPRPZkNpJEqfnb4BpUODpgPfBsprmYh5zL9wDQ1o5dHJ09dmwsjL7zt1Yu
TNQQPA/pbVUPsPh/sKq+/qXY56GGbTGGfKThbdbz0A7IWmjNhvkvEJdf1VZ047GB
YdE/V6vSSsaz8CjascoNcRr/2VA/9kqJRqi3vgbtgrl+tQdR0+aKSfRzIENeYeQl
3wcueK8TejJUC/fpZGgGP6K952q4Di8d1FXR5BJPdMJilcZiMaMSvR6Dn/oN5icM
rytUChx/vQsmdsSCX2Z/ykKGbIC2+Qzm8t1ZK9WawrUiM1gGghrsNM4nJTyoRK9Z
FoEuknYMz2NVsU3hIuX4qFsAawmYGW/B3P/7HEzB9aEVpfAe6693obZkRiupYnvF
3hoNYfkRhDxF9u0HxIyUZTWAJ11LhrSAPV1ibW8qxtrxKF7pXirc6RzVAyjn2kDx
DPmwmD5Os0vRbzlUCFbQK9zRBjWe35q8xapuvczrexx+AWA6QdNSoywEh/RaSY+l
veIHVYPLNvl6fpj22pqsS8QmYarQbxxusxJWEtpLtzSkGbsjQlUlu4CtlWjUmWwl
YvPB3bLk2vPF+E2+N+NrKN8iPqZmcRJEKbsPBrBGOD5XgIEG3sHPed+DduYGzb99
JL40+wCadwMLSCqeJnFY/pwcDB7/ALBwYRraVM1LRwJCAFI6THTma7HMPM1j7C7e
1dhYB8QF/Y+pRtHRterksLf0cBC9QVvi1K6biNlvKx0zQcKtj+ywPpUlZuG/1iAN
eywqUIplavjOAKS0DfFGI6X5FOtO4VNMLlAO0T+nZiwFEifW6fqzg2GsixRBvmxa
/3zpW59QGG1oIk/gjeOcG5l/yEr344FKoHHuhmAd55BkvAAjihAAJlwKHDlXshhU
hu3ZSUn4ZzA66hwWdnFXXv/sXgXIL2n5yua4jY9cUZ0u/3pBjQ8mgV/uFSQUKeDs
3cH1L0jxkP2Cm3ihQgk5jfu68LzjHiKBNWcvAKVU4sgfEnfVNAMzrJd58Nyu5t7H
3/g2U6EiAJGtJ1JU4C456poA8AZYwa1BZFO0zl/CuAd6frcSdh2evHZXJtCSP47e
/GZymxbOPrSJ5WKPdUs7xC/Zh/rH1mgeD9lbgYqB3T6Uszbw6f0YbweOZO5+xFc9
CSOwm+m7j3Gm+cX5o7W3MrFONBxVqEFWe8JLUMMY8Jx3opeFrSSl7mDcDLGoGv3f
lF83U73LBosKKvuXvQJbebDKm1n/Nxdf+wQiYafXP2eCN3nt0tb4L7x8xEJOhWgg
dYQaxyuddDJqjn3lpteq0Nvq8gUBSJLvYju1leTKdBR6RlxPR1r2M4RdjFyy66AB
tQ2B+W2D66qkImczSe8kcEvAi9Kwj42slxehlJqSlueI39s3N8zB8u+sIYvOQBZZ
2N8KZp960xLXs+1R7EYFTdOaU35f9wDtP+mqis6zoKDm/up4EuzOvRsmcuKNPV+H
ArTIogdntjVzIQzHNrKx2BF6TDWV/hSrtIyCFlkKagaaf/WoOzWVjFezKQ9evM6U
zpaPg98NDqgfCHHzzHLmKZDv6PYpc82zqza+/0OsGWLsEkz47/lrEs64La2QJpDn
GoEdAs92TqctyNAJirVRqV7N29hhdxiyVLuA72DTskD9mIbMRCX6S8hk9iAhk/i9
/fKicsYPnt2FhX1TYMTWVR845iZr6X+S1F2W2a1Bt9tCE2/kUKnBJLZlqk9XaIlc
YfDPPneyQJYnPXrH4hJqfXZOP1kjZw4zSW7K2nzhhve05hJavesZ7aX5FsSrPNIh
Jwv5riY8ZlwA355mGYZxyuHJmj5ed5gg5pG53xY05V85RgN6p6xInqhl9bQnkv+i
h81SovmyBjoUp2k903pfRHYUWAl00CHIqEiz5vwHp7BJgDS9jwAJM+Ke9l2mvoiN
Qeb9ZqUH7pWGnCuo4cBFm/Cb6Ktwr/Pt3CWHY9FcQwMk4C7KbAKMTk12Qll3LkkQ
NwvFEvx1RezeqbT0C6U1O+l8WIiBlLvS9xaCyxyVu545zvFSlITf571aL4eXRtWW
P4CWpDBuXrr/fK9cX3E/8aZ3Zxzpn06XLvmsvoQZdq+O3TTm5oJPwE/+jX60y0HB
Ui9excKOnYdx6mgdlvDPQUWVg7288BrXmzzsgGdVN9Wwx0x89XDa5znCOjnPbIZj
NwfE1lKbSeZ4ixnRT24PXMIJwyyws7nmJo5EC0q0p61kFqgZkvLt0QWAEy8JdwwW
Ti5yvVmac1nzbQu5+7+/4+1r8YVi5Ca2E1z9o/eaAwP9ivh1UDiU23w/hTaVJFk3
NACm+KTndGqT2r85FNxtTv0p0Yq0lgyaPRrCdElmjB2mR8Xe3olwGrzZiq/u86DY
r/Yx4yCnj0dxf8hwx7FS2/h1kWsjCLdXal91LQazB27dhBqcWHMdcLA0F5eLdEmJ
rqi1hf5ZBg4PAivGW0FhwC7PhShSoTmKXVEq007c5maVKwbb2Hkude1ZwKsw6XD2
b7oLgnTl9b9GZbEVredePz38aIzdwx8pJAzl0EWrUpMwtCPTpegpjE11HQqs4RbW
sAypM/mBGXwN7Hyd7H+gQOAcbiftTDUb+jbR3LsmikL760SnnjJJyI8FCWVki2UZ
uoxkNuy2FInGN1JXxE7Rb35rCKgOf6dlJxGxlS6weRRwEaR/gULgi27rJl2hXD+I
LqB3QxasuqMhhdk4JZiN1nRI/3zUmk0JAN7eR7AP6DHDSWyQcRNuLwBZ1DqVNZ2y
ZPwGVJx1h2ifWK2osSiA4uk84VAZyrAI4jcZ+y3EGU/HahjioDqo98+tN2EaTWDk
3TfVef5hX9/HjkH3wlz5EH2tUkASxJJikz2phQDHAVbWNBOFlzZeF7dupK7PhOFE
eU61kaFnBN1rMHTFK1b/XNhzWNbUabTV40j0tboUBRw6LL160jEoXQeIEVwTiEup
PvXNQLuIqTAwW6/uEo8K030IDh0s6vrswtcqToGTVZU/C2jXjAp7J+VdFjmuKOGx
oiIg+Hz4u6yqhLVNymXG00EVyOkS/KTfzqWdeQYaFA+poykjAvWLinP9Q/J3pUGL
uIQ+qIED0sDIr3eYvJNKlHgAFtEwPZHTRrbhFFLZ1b2crjWUdNl8BqB6AuXOQd2s
f8JPJz7a7VkMYfFS9a0II6cxasG8oNThvy2x4VKZRaGBo5MvZNwb7m/eq2x+Thr/
moyVBYTRbvcey/AEutEefPBBSwJtay1Za0DxQXrzpaBokJ6m6zZDRqElqmysNplR
i5XKW5tLds7XxRHMyEMzonz0V9G3ZpvikvB14SFFlycfoW65ygVraoiqB5bNFNoY
o0suXx6NsjqoR0jTBuOK/hXWpPLmTbB+aId9L0rt+/Cl9SuEmzFCdEQJaroAVqa2
9i+lDw1IrS6zQB60kiM5zilROVekaSNHZ7xq/xZiCeOsxTQj74aMxAKisZNF0yFc
zSj/MlNoxmFY2O2WnLPkGpZxGpC17hCqo7PkARAQW/pcim/1G53VsBC17IC0c3d4
PlDO6bcAyPRLnSRx4lk2RphDX/RhnXR0xtWt1fDVwSYwlaGXGXYu/OJwwqfhSzrV
sxenA0jh00fy7cBHejY49zBzKluMEhQVeoOUMD+fjz5IQLHhHPEtnq+5CcyXoL4A
eYT+JRZq1Q9meBuPzq+Juibi0YSLpqtBpJwTIfM6JCMOr1tjsa7Dsym3hV6AE1X4
jyTv3qBSr4+0KnI6wAwXm/tNQfbh1DH7XiklyXHRydE7jdaFdVY3dnElGha2YT8N
95d3KtcZ0EvnqGrNbKcx/2rtXnvgeJzL6DgrGVumtKfVs7j5kWBzKzaWsNr1CdQl
oTw/Np2P9o56+nEk67gML+EuBfhBI9XakvoKRXPki21r+b14r8YuNbl+DYd1aOFt
cyNIjFklv+qPUDzvckSbCCEAAi6O31a+qpne2/72HhXd+GjEktDgg5mK0rKIRIhh
Dn7kmL8y3hyPr+yiFVxVHCUIIR/lmvN43Yc+DKlAn5VSZK1vPpWi1d1498E1FMSG
KzqNIBgXtnxFRffljiPhA+5BUEyKZpumTOmL0Toih77nKKCdQ2IXSwXUTN5tjOsB
eDBJr5OWXWUEbK0Ay+X5SpsaPWyWd80b2NR6ZvppWFK12pJ1UqT//hZ7z5iMpw6b
eW+OYOVnKO3NbQghcVf7vci8s6osvC6vtVigRZp0iEM9AQYN2RGeUMBBrcIY7KSx
T/zsidT5SAZDu/mbyB4l/fZQjmsG/LWhlQ1IaDgpk576zGVfXgLfjWWUol4wqHHU
aHflTd56tOTc25Zo17tCZ8Q6V9XqVepzm3tPVO7FHe3Otvw/X4CIotkhRhbGJS10
1tiRdKpfJbkZtg7eK1A222dU79GCwpWNvmGH2B6hG2FK4HJz1CkpHcszirJV5+T3
utQX9n/Za+ad7B4aNYLWf8yqrHfOVXD8AzuFzOlmcw0Bg2gGu37AgD7doiY58GKe
GUxr3vCTILG4pu6UxWLDEEGbEEExuCYYmeKwlWevcP2Obt3IXC/dvcE1TLFT3SDE
WOD3pBYFMLQjUSnfkQ05/1R1F7MhTzEtmEjEre9v/RAwmfAHDbdHdjWsreC4d+7A
7XlQoHFqBnOU6ppORY8VySvpvZuBdeeU3gMNBeD6laKV1Vzan8+5lLi3K7kxrzE8
gANeZxFATze6Q5wg3zeKPrtta+teFH5tdh9B+bYN+hio44PBKV3GhBKCLCNEFb0X
9YWMyB/RTKH37gI6RRuzhNik7MKBUfmmWJgsuN07tC0XQJDN4be2BhS9hKLkYRgx
RZ1gEadaAtDEP3KuZh6dBkBRtJpO+kq+5RzRvysRhBzaNILjalcsZWAp9r2ak/Ds
RGjyUruoDWGByn0eLtE7moGOLz6kbMSMfVFoqM5sAm8A9qQOGTTfMuOQnjNkygHZ
9ZYPjGrPO+5xxJA5XMNcgJQpPRMBJZQkFqSaw/l5hsGH/eKtUfNTf5N0S7Hozy8h
nND74jV+OSttYZGRoNPLszidjN0Qq3mZhqUFLTMSwJyo80siyYFxw3kzYxVoIXSx
m0PJyhcddLwWTNR0YlD2UVcb4MOuZa4tCzESlHt21U4NebSrIKi1WXQZNvUtY4t7
Qzx7IdpkTHpPZ/R3MkKLg97/3Z9LdKrsOMBRn3z0g19msn26DPx9tHYjntTE0rE4
3MwiTdamnqSEuJyWm9d6RCTyD+CRPh2zX/F37MrU+EMcG6IgYyGVa3KOP15SjQHU
YLoeQwSTl9Rt/nJllf8pIkenc0125TGF3s6up9fmNP1/WO85lP/bhD3M5ypFNQZ6
4PeNVPLnzPVGAP/eTdlIqkuGuLrgei2AtMjFNxURmc4pySgjNuy9nJjjgCH7yUCz
6H/WdX9Lyamt4qdxnlYzkfaWMV7XcIEVoGrWez43oPrjDfVv0zZhQq7BeKsRFMpR
B2v5FTB/L1d0WOlO3XP4b2CBco7M2af2TrAElOIxN988An8WhdNGqIQAAhcjdu98
yN68GiwFdBbPbdQLTB+SR6TAwv5jOHbBQ3/4Ng0/Uhi1myUrXvUKNWIVMki8X7tp
poRFUlkTkRZH/Lxs7Y1gizWRm4TcuwjEP5t7CHJtNuoOfE7EnevAklVnWXQRFt1Z
g20yoNlnFk6lahEWKUEXr6el0VVwHxMeNElNVrm/rU5Ruzr5sFa9lrrjWifzCVJk
dEozz2JxiwNvUeK/AEmmJFiKdfykQWr7bVm6n+F4WBdrDtSLczlASXUCqtyXty8z
/M6NDOaDi5yZ53tBDlsEk0tUx12xzebXd6a0ayIUYD0jNvZPEdb3txsKkZP3LPGU
Xq+aBOEFArpdyD5uUpNDUYVqlqN9bQviArH699Eth28UAuPiJj9KQBgs4SIN5q5O
vfOa5V1irH4zSjSKXxNe8FaleBgs0YdSkA1zAg+rQNp0rc6I7WiHT9wgelJK2ujy
dSfyUoTG1rY1Ces1QGz2H0+mG+2r9UMD1i2wJXIYWkqGAoJgKAXfovsIsQ1LH+PM
lk3bZ4uJnTlowB+m9ZM2bfRFoUtkb0cZb9kFNDtDNMH+rTPqhJ8TqjeQDxXWS4w/
+27MxEKb8XVcVjyaZVdw/4ejnFKfc7rIWF/urYR20Y01mi9Je0bgThXgEGKVIPLH
BLYO4EAv3sRd6MaIIK3TjzNIQz0A5s0D8xYs5PC0OceflxakpxqEsRGncctNWdtZ
uUmmhys4pXnO9Iw4UD3BMalxqTizNE1ElhWNkXS52/1ylqzMOgyyjNtL7Hmvo5xm
MiTiiJA1xD/hoMzIg8v9G6DxxC59t3HgB8H0o4PZQmSAYMY22WfyMkXsF/F/atZq
iAJFrVmK6NRlfTDMBB10TMscc3zycKfIMasUTRxeiemFgmOv6Y+7inBx701FaP72
05M07UsH3UoFCSzwaspYeZkNFK1/F83BTlIlduYLDYrrLxaFGH5emdiWgPCZ/slc
6QYOWhe4T1+n2xGZvyBCJvuWhr4Pw2LNmC4E3V56Soob2M9fnDwI41QRlJwNIfrP
43GOFPIhsHWNrJqgu2awNnfiIVIto5wjNNWEMlDACivXZpbkfNMH7XPbnbUcpeEY
KA8zDBinDX2ZYNXKM/+4jlxlDd6IMxL7QEZ5LGLWyw88RO09oBzS5XJhPL9bSOQq
ph95M/6OoQZ0AbJ9c35afTUKz93rjaAjyl2htF3lEeKNQNQ7rvputW4/3MfeSCfv
xUctJ923I6uy6zzkOifXY5Pj+OvgaM/vTlpEb+7e67y8/5dNo4eNATTkqZjW2vtl
nSssq/0F2LwxRYPor7zr0F2iG+/LjBHx5HwrBu7fKZfx3K0yRx5lFld0hfMQXCes
PJtaCHddzqfW0tFNYiSx2g+eXV36//24cgT2/GTDn20DKy3AqkDxvTUfZO3Ppo3h
/ZWTVj2Bwv0cb2bfqXO2dHJLVAb7xLhq3jhFF4fNdOkzZa0mm2e+aGknwz/IgI+4
Cob6ccGKffjR6ujXJdnl7H8YjmDnrYAmDZf9mCpJLk0xcu2ZFcUVjWjw9Bfad+VO
mnqxtXDqv6kcMuUwSHaLJ49B0xwhhptZE7FtSD8Zaws27jvCO0ydZHAZ4p71gJod
MkfnLMIhV5ZIeU5uNHTnblIE5UkB+t7YwbSuETJJyHPrV8udIPlWZdpOWlGYl5LJ
ojm4rmiUJMldnXbpZVky660iKSyFtiNXNLZewCeBGuH6bn8UHv6BKRCVwmzdubDv
wHl7ElyEgrnVwZGB9675avQkOKCdQ2cbpNJKWgsVV7xTfXgyDOgrhDglUT4t2QzZ
Nxyvo3XDjnTQqijxcM4hobJgNnBBP5rBesRDzCnK58e7gFqrO0jib2b7WYbli5iL
IwhSFwvkL/QtXbEBAZb9wRhePMxm1qh7UID1LiVES7LfmVjIoMYn8MjRLq4VjYL+
LgGHuQH2+1f8heegobStkbLjJmAWTF7GdGSl1rXkrk2joi6xqfVxTARQR0nKflw2
8DBBGaZ0lzCvY/+bjbjo0abNgvbt4ZrFR/VCJvIO+31Fn3FF5Y9T/OL2st4Ganij
pqXN71wnCHfzD5+Kdd/fnMihEGmJBo6zAPP9zlUyhEN9Pn7SdhRCimrYikICWD51
iD6ZHp2QEul1+R/JvdXck0WB8POQHmBF4oyD267gSWzEJ0qPyCRAb44w3uDkEVDn
hXPlaTRSqbap2vdnZo26n1PhlHF5LExoxVFdYRHLa6TfvAkpm3H4CZkG5Avpqco2
m8c5utX2pO6Nd2m3hTgf2+ovMtggSsZoVLmrQJA+UGAfrXSk2OlhEXfNXd0QWxnw
+5XSh8QUX8q/+xYfwrWtk0OJG0UUszt6dEPlP8649dY97t3HoIMq0vrhL+VAePzb
si93A/y+/BkaZjDl5lnBOPPz6ncBPEoKodATxc0hVt6SOORD6Wm1LU1j6NXs8TFn
WoSQV7HBXwCpU2W6bNFLAr9Q9WppvDf1q63TMq2v/JiJfOg7SfT5tJwvgmwMMKvK
4rCl2Pq09FYVlcjaX+6bz4lkulUGTyXAOapwU5NOhrQIC5LDVdKF4v5o0uPepB99
CC9Q1Kf7sYp7Wx/tzONe9gbZg6gYGy1wM3FEtDdK82oDt/hP3UUDrFExYGDNcqKM
HbcvvFN1hCPSEx3FSxatupZwcnKgITn6c7s/LBdJZ0/jPegS3r3YikhHZWFgWy2k
4YpfkQD5J5pWDZAGSGE3rJXgtnMZF1huXkWbIBVmR243Vh2asJs5N4l3AoHh+7wI
LGhMEJD4lRztIrASqcnjy2g6nsDsqv1B93OV2Dri+PtuDnKJ+NTEpKb5RJvs+drL
JwZy0ZzKR4baIqkFMny5sCQwL/5qOhyYEp2VbMO/P3M0fU0DSPuuPAWEh1goLpjm
bfnuCdfPeQVWOHwWWGpd9Z3RQjMd1c2tUScDnbdIlr0jrJ8HvpTTtkMJxdQUFhMe
yOTyO1QmLpTlZ2ZLX3+XBoZC1Q5Xumyr/MpwDeEj82+clyA7Kjmdg0ednjpA33W0
6Jpez051//QhkmMGnFS9iR8LqGXYSKLjr4lDsIHkYjPXbfgrELT1zZYnvK9PQgqF
OaRFb71E9GK76GcItq8lAxdB/tJHJzrysgN8xg7kR5DSYspiCJJ0F+bkQjxAbEXM
pNp7CTyw0JELCxzd9WTqWFhsXpuITsl5wuA1OCwgAHw9CdO95qGdx+2h4jiK67RQ
gY62oucvyicAJ8YvJc/p3g4wFvnF5CEH2kJzd/ooEbu81GQHVUb4+t0G/xmuW3Cj
wANye2bv/mdyktTuOK8/NKs03eWdPdZcqa4t8I6rb+4PCK00/QghJ5e4DeNM5fTA
Ab1FT3IkbWSc1hCKbkl3KpCTqbohAAl5T0S13tk2am6Bo8TxMX64Vhn6uTCm2HR4
D6DkmIoq+3BFGUtoGE+6XrtdbfpUZPJM55gwl7uKle6PZEORguZA8LIdv4bx+WaX
7Me8Gfie8Z1CSvHADc0bKh/JwLeA+q7VcGKQDgsvmzfWC8/XAcLMY2tlu+nxZ8zm
Z57C3pyA2gsys3eJnEfO/NCTvzZ/CberuhtoCwORqTxWqWKDXfCdr68HGDtbesyn
c/KU2nSxVpu+I51brJoo77G08AWFMy1ecsrQtSuwTqJRH6kdn4n+rZw+O4JOdM5I
17PJs5tUJ/A3YQ2K9WN/0REVAtqTrRhupZarht/I2zR45M/x+bq08aW9ejQUeoZn
ncRndhamWvgLDPw5Sz+59Z3Djq7RlqSPAjDlJ1XNQeZ7Z4nl+qCRbUwXVd3LRsZZ
dBiPWrfjJy7K+RVyQEyKOXDKcLQPlk2MeSa3HMIrtIbppjur/KzQ9XgHZVgbIvB0
rgxQctyt1dHdhGfHBU7APJE8gQbatPX2ELClle6pEMLw3RvIVqOOzNBENFQWwd5K
pHL2hRFqZzihFyT4N100CzzXzU7vrGoJZEwg+FID0yNkOcgxs6fOaJismi/h7H6H
IqVRMtYvrR76gxB+mgCGdR5+ZpF01pM8r1AMPRIdlZCDBUcF4aM83GfjGtzg7X3N
hx/Lbyx4CS2BH5neCejQOkrTv78vd8NO9sSEtEypacQMlijyDM0HiMXADI/4vwa/
mlb1SROMOxWrMn1p0FCBqWtYbR/mkPtvHT3sWiC5igzrDsNpRj4N4Vkw5EgexkYH
HU93cd8RWiuD0nrYDunIyob0mznfi2Stlq2oQWlq7g7jrxd1QAEq5+oxIUR8fVtv
4QKmv0Ce/llqKAjs9YnoByFd8yqGxdMVE/eblbFfE29vknKTqgxUQ5sqOi/fQROd
EqhiKKtcARpU6Erhd0YgVVAc2tpPiQxts2Gf7+9A24coe1Z1NVX4LYSjBqI6RQnW
lpddmmmBcJ+jZBQPe7tJLSgwbrLJGvHFyQMKAxYPsI8jNKHwVulhmRj/6sK3SEbU
xsbXZzrauqkS8hRJsSRfJF6KVu0Br6d0oRCGzIJ2ksgCj+pD86KWDQ1ctC0q1Url
Gf9yvOVikSMSuG0PIZ9W8Gm9B1q/qWnIBfkRJT6j9powdVchJuKprt8/Wukm3wJt
iS1ab9GaqaxUYHnwaT2FhBAJAfSSUW76uIKSfVEj10676m3ZcC90Ni8l9Tzby4UQ
xV12sP4caNTkydCMT04PPWZ5X9zQb4UU/ERIzTwqei2aK8FQyT3rrbUfCn8GL3Z7
aJ7iaDovPThvKc8+NqBKCLP6NsaLYE6Dj/5uGRS6tWxQniUCNflS6HizI2dKQJ3Z
8qw79N1uMt+mgIE5kEXtrffFf4Fva9S7DoSpbbhxT0rOqqh0eaPbERoBXze5OHeS
ohuZdCwuZGwpUZeZOjfDQo60wBZK7Zh1fQBonUox+n2slbjhk0rApq8x2MA05wU6
fu+/HWQCLbkcTzLq4lCdbYkssGIdDepFc+fRi6IwE88F4J6AnDDHxZQ30hKbb2KW
uhZu4WRkPrgVCtSm/D+xiGwnb5LDBq6NHSjMhHhbqL9FOUWvAhBNk4PLkc+7H8wN
8gH/xNvDf0R53VeKHZV2YMwG6ry1zeieXpc3MD2FCoxz++7r87LvvyzLOxkcpRha
pQ5J8iQR/tsm4AU+S8TZITjnIKMleJgjNzhboY9SZeJ6CL0ltFnO5mgggMr+S6Nw
qKuvjdlmWPtpxg+8T37CijrngoAly/OfOpEaIxsZoTZp3jf4AWaTDqmfo4t37SuF
1MXA6t6peast6bZaXWCUb0Ms40IfO/2h257zRYMrPeT7glazDiDiEDFOPFReuYpB
QggSahjPlYADDjhy293cET7Y4oOgVSBE8IrXYqIlEmXrJbkHivX6WvS0b1xEHdU8
p06gnpSZLYy8Af3yAwGAh0wq3D4GK4Ki/sbRZYhbe3/eimukfDcANHqGvP2n73O+
tmeoNmdwBOF1nKdwOqhYhtoWkN09C3P4pT0T0JeQrOw3ddFHCn34GPh6T6x9x/V6
ETXDvbBhbYTBTck371L50hI/aZPRe3h9t1PI4m0p6kYuZi/PK/OhreIMy+umkTgR
/4TnUadE1ArmaJWbLkWwJ3WUPNhdblw0MlOGzxO7RYu+v0g3st43DBio1nqGmGRH
v3EWQgUvEdm10F5MCHi1jclTS3hxz/c5gMk3eEOwTuBtuO9ipyUN+gZu+KWHtUBn
pXWuG7nzgiG1x1pdih0YhFQK72ZZF0W4IhORvB/++KrxRJdVFfTjSV0Ck5yobpa2
M0yjzwe8XjWeZdtDhcwOx0Qamtl9nDKfWxHbly70mL7hJ+67FvCz8IlUHAl6lZRt
03tMcsiHeCxuLwM+6xdz7Fk9pX0sJrtY7QN105HH3+he0WzMn4RMRdq4TwC47N2j
NezU3uP+a21S3Rd3m3ySVuPU+CxNkG4HgWwB4OniSYxPJvA14JUEGKxzIFBTBIwe
75+cv6lD8TQkNvEBCnmQRVLm4okJYbOFxQKaRRihf2Czfh8XrZSLFP5aOW3LMUpW
7b4aeLbElUE5lL1auCPQXt5mUFLWu+e4EqwReE7oaiXYv0gyAmaFdeVVJk/9cVMK
m2jXye3dtIzHplNryWy7q0gkNFBch5zEwE90oCHpF4R1J/YnjWjmQF6JHvBQ62rX
UV3ARcSXAhkwa1uaDDN82kPqUi+cqeMQiNu6f8dODXpr+9AEnwm0sPGyW84QFsiS
Cv67AqkTh2m4MJSSRS5vvu46vHc1ph1aIyBgrONj/lY8LRPqTpPSt9ncpGcYgdAH
MhctHCP1k0nTYJIBMoAIKewHFhWFE+KvUfc/BCic+HogTz2w/2p6paGdc7Q8tEu4
AcYgTIr5bsK5XfyOeuB2PJRnEKjMpXgqC+qWTNJ6A3/V+a8SJe2CrDAJ52yEnui7
2CP+TTQX2rJwcLzyr/hpH+a32D2+E7T/9ZgWvmFczxUAeO3BQSW1Hi1P0/jTNiWI
nAhTxAW/FuGX1Zi61MS68O4YkFkS6nsGzsZZZsxgk+qavq45gw/WW85tU1bUoYX4
peCeqfpX/jJqcaeL1biv+Wdv0KGOswYsTPFDHeZ542+iFuM3CY8nSCdlnZ7Kb8+g
CBsyLL4p+x9D6ABA+Sfth5xQMMGDhrwgPP3VGo/vI8XTeExnxhIIEC1RJeSAnR+G
54kP029jsT/P9rfGS4GnM/HigATwB1vNyb++c1U83WzVdC4gDKBe2RjX5hGOppFv
LWj7/Fc46uN+HssbNPju9g7ETjNAJsKcV7JBdGlVQpmjUZGcBsei92KJTQgSg9As
v+Iah7e3LYttlultIu1AJ49HpBeNkEziOj1fQ+WSDOsEf6zfI9NktUhroSSg5UTn
EdWo8+usmlGaoa2SXbsavzlfG60Pf6UjlwoaOBGIpCM1XfMF2Z0bHzyv8bKjCm1b
rWMaRoeFKoknL+GlMGPv4wlLnTuNjetK2uydmw0qW6w7OHKjDG/WI9h6pcJuh/2o
Dz+k/6Lk6EXJMAJbIaxVOFez50S3bDo4j+yE07H1lTT6Nek22lRzxUG9YilowyNU
+0qXVIhL2ecfbgbOyJbEIRSAnsXFSpkByfRNGbAEuX+oqiGruLArvgqj680DaB+G
7dDKBPViytVLs6rRp43MhizGqF67m0DYF5lfAGZd53uukWnJrcO67AHBbKR9HsjR
JdSVeyBc0bjKrM+dgcUOnXcbPH7vDJrAtXSR3WxjD1Xrtvp2fy8hrHM0Zw+267RW
cXq8B1gi90rNwcZx52A1Bvj74vJtQ+G23UBQzFRF4kSn19zKw0DeZOoMIIiEpkZP
9ii4ob4FmmxGkG5gS8odCtoPmH3FBkh1SvrHQ+uXor36xi8uM7Z1NjnDxzS1MLO0
T02ZCcpe+7eJphyIZk2oSws3Oi90M1Or00pgtY4zrpqyLPQCk/hUlIKR9vKfL/E9
1a1ERR+2zZAUEp31Gz+Agou1VIZ7Nji9Nf12uzDdgqRc5acQM5iKSQwhZuB5RJoV
lz/QoplRysClF0uPxL+GqOGCRdykTQ3xInCUjPC4XF/GUodRS0hin35QeK9zm4is
YmvjlUziSQQa57XlC+I9+zAHTq95qCm6TgTfuRfBmolScmSMJx4agztRZyWa3/X4
bzZ2yBXmw2ZVxSz5KwtQMt2mTVIyyzQWNxFDstUwDyoGs8Bin45lOYNU9RvKiyTg
Qa5w2mzV9W5apugBTngGf1rRVS3O9iQO3LsoOvtkdo2jdiED2HlN7nqkIic7yxdO
Yy1w9fw+UBOF2slL2uln1QPSUkdbiXQeuZyKVkC0kKCoLS98vg8/UaNaXTnSTHUI
/6GDMmt2e3anDnPN2LVzgzEhNnxAlduuarsqtO4MAnBSK1V5CCidyXuHPqpAPCTT
3FpMWihmifW2TfIxsi49C8mbZVMeLiAkk+nV3B0ufk4TpAq4sHzBzU+oFp/ossDx
t6GAbjwFkT643GhSCW7+VDieRHcKxH1lrJ26WhbaNDRS20mtEQ04GzF0Eodngys6
T8Rvl3yYErSOsBXC1gpH088/yClmmFa13gk8FnPVyeuO47r0utdgGFRXRgeQC9y1
n7gdEkNF7mQ9zK082XYIyxS6IlHU+B+Jbw7srsfbWgiitXw05PcBVi6n2cqJx5TF
kfA0HGRA/i5YRD2fENEWLz1IJrg1jn18ULoPRybU423t+C073nfWH+E1jnekwa9c
8BQRLrgulw9kvCgFL9D0vQEwlqXqaCVPl8NGEsv4HzQ1BhOttRLnFFESa8antiUY
FwcGZgKfzeCREfBmRF3+VfQx4y2Vk07CZ38J6Zx7iVRzapyH1GPaDIXwVjw6CkZE
henp1RW1WpHfm+ZIneIO8IDeShBgbQX8Lof77oGioQykv+0njWING5QifOPE2HbJ
w+e0JHRuYqPj58yEKUBJKjmMip1ovlZEKsHQFHRiZvUFZuKwgZLZwkHAcU3ItgyR
tUy0EBf5af3O9XWaxN8hiQZjTnHWEhrABaKmeHqqZHxncXN9efa0cS+Vbn3FGxaI
Nj6JOtOKjfSxA7e5vkKVvnz7E/gUN4A/QViA+EIfQKyCEcG3qiDmP0aeeZb9jGyY
yIzaYcMS6PTYrICmsyQe6lpQzJqMvoYiRFWVleIHnMNdEAbZjP4Exg1XdrgeDXcy
JDhyqp4CHgYBJy748SxBEtcWWApeTptdNnrSLzhTMTaXU2TB++nL+sE3gK7J1wRK
RNe3gtzSio3SH8tCYlZ8HcpUvMapyT89AC0068otdnmLn/wAzMNmVy4sFbEQuSkQ
AmsBHGQdhNpRSTOLOWYKQcoggv5sTgKMHL9kzX+f6HqFCk03BcTndJwMNrcLQvKQ
Yuw5urT76Wm+qJHkqczi4CgNGOj0l++/MiPzwg0D8ui/9Q6jBE8vQG8MpvOJdGh6
t3d4obYFtY8VGPxcVPdOYSY3exNqnAQTwreyT560GFK14hN1A00/UYWTGyEnMduQ
02QVSp91/Tve9vxoFpI6BAFQr6aX9YIh8BSEfvyUnR4O5aZUFcmukyUsEhEf1A1X
kHYmEadyf/vQDZwjIk+aNpqCeJi1jTdBUEg0WGjYQS4YFKWz9hSnSfquZ8uzorXm
YwS0eNBMOlqRglirSH3B8wKWypexfdui6EVlLsdblVRIah00Vtl9XIhWKUS81xtz
uAjknsUm3wSr1h6uUJhuLghiPl+bTLyi+0mvxLEOoTOG9fessviq3/TLyeYag0Ef
AN1EsT5e2DGa2sKcDguG8I8JViO9MXsdofit+V6kH7PFfe85Ia7p6ccpZFnCLCEO
x7kzuaEaT4nEzJ6OWsFSrS/qr4wLpfUl6vjNtHMwCy2GUiNeuKiBDbo2uYiApsom
0AgkgHGAh5iMiSKMIQ4aeRuHpO6sTncfdXb9fHl+Mo4xQQVfBU49+1+7grHMa/XA
nJUgQ8vg4cQeUi13UanXYnRCR1G636bTzudBcYm0F9itPgsDkSjV135P/OKX/SkZ
dGj1f/3vVFmaIAcX5yqx2m1KEHdStrx2AFzJ80CNP/zj94hCY0RjB60Ug3z1aCli
DOgOErm/+qF12ysLVdAj+a6OcsFaLllEYgtkf2/9+jX0uYIZmVCuzWAaUkVlsuEs
Klz+hnlGM/1GrYviY8F2UjLq/aYqQAxnvP+7JEmPcMLz160oQjARJHxDAiSm5OUb
2483zXwe7gcXqOpmbnRhVbu1yNYQIrvgd+5AOs8iFQG3Nza7i3m4cGTIUGJVJqp8
P6HgsoCK0X6YrYyRSvnw1pyckOKuYAbCajHshxZQXPzUNI24PccPbSCs5BZ7WQUm
Rp8De9cEUhd/xEWQYfDDSIa98oonXxqz0BZc0xIN3TBf6jDy39snywK0m9b71ult
u2wkhjAIEkib4bx83yqXL0LqT3DTpj7zi5/Oz+5CLOzsJxtYPdHZQQOr6/5oam1q
OGMrRtnHk/RdimiwpA92VHnP65tMTb1/7Gz5lT3P7gxIFHhOtvN3S+iTrYKpSFUX
7xAB6UynOiXw5iR+1E5lTv9ijhLZuVL7k556mmmdjkPkmZd8/F9ujZfR73zMMVzw
OgZYOeFxA1/28q9fmNPGb6onqkMKfQRzGdcZerbhBFNipj0z5bPQMfL0e6oMPzMb
kSk/4bf+KYByabeQef+WIUrb0x1ojJw6uY1g3TTNx0uwGH/s9n1GbAichx8To/i4
ndlMq0iTIiKhtU+v9qeOKr+ZC5eQcOGaozpVPThE+pHE13UmY6ZjtACP5z8Dxee3
53pL/cmsu1CUiflqEURICOHKxtUoyZQ84a3uTiDQ/gYtWsMCqYPD9FUixyINdELt
+iK1yajNYZxtMgKNnHMy86VUsTBSzZax2QBKzWPovzMVXBRg8hG2fnPVmQr/YzcG
dj28ucI5+JCoX4yffp1UXpRTPejqIGuwHqO/flQ2jkII3Cfg8+skVxcJLnHxGrWl
I9M2seq8GT+M0+KHEuifKXh5fd/NpAkUEdJSuBBbRieLFbDliq1g4Y4saFQvvqzj
5TCBL1iT0xOavvCvliMxc6LQd2ZJCDEnwOe2ETL+K3cQyxt/WayyHOLCt+meYc5w
tTKMSTkddozGp8ksVBPW+9uuf+pKYNFbpV6zhkT1+X4NZOq3iUutgr9ZWtJZYJOO
pfU59UwLyuqUtsRNTvn2lGxlHLhOmdGBUshc0Xf+4NsPPdLWRFXTAWXD7ZCyRu8k
ZIU/1ebTG85YA0R5p6nq41M8Rosumu+ruufjoaASsDs0qKiVvOV0L2QTVBPer2yc
XNKsve9GxnnTlRk4eBq4un4fKIuSoRNQakud8o3LqJpYJ7sVEAX2qQBAcI3estoa
4+Rd1N0K2Dr4Mw3JQxA1UnePH8eMOKrAVRwvTBKxCsqS/IVT0OCKyOppIW8+Y5oC
xW9C1Ccj0sLSA2AavZ+VdUaG7f/gkiFiW7evdOCUjimFmA41TIhae3WU2/nihezI
4Idhi0M5OX27YEn53ksHkeFqZKIHpwsyPcJvHwjlXiFPWrZYFk9klKYQ5JI86NgW
F6GoLfQESoeD6EnvoFgISm9mwj5e9JMDhSmJk+Tmb8SmD24OhZnuUeXXjd3fpN9A
2vixvsXJFc0crb9iFBWzmveLL0ndMVHpH/yJ3m8rizuf9LgBTeaqGSLngbQ4LcKz
Kf221sntktMRwzQltTNd5sI5a136ZUI1oMTla/DN7ME2kMo7q9vreB9MSe+dGeli
hHN3QM4mX2xr2MaYpLNfQKXkDWCLbAwDqA8pdcyg4zLYhtFvDkboSjnU2GgJ7FCC
wCIMAGG83KqmAJ2abgdHa5xKBBi5EmE5BBNqCHzGNBlDHj9D77RqDv1KUmbEBxWJ
IOyi6eRK7BAwNM61it4bvWWxBodEaWih4VS2ifyynfPAtRsAt7NY3yQcQO3/EzHv
3Yg22mwQNFKmjkMAzO5TnzOQ2Ipp40sD+RvHlFTdAq+/tRmnJmxzG4dMKlaq/HcG
JhXJMYmp92pdyACmyECsQpOJVpH88Ou9em/AJCesY1Eq4FLYk0nU5+QdfUX3DUSv
ZjpVufXygNXPc7svQ8C5dN0l5StM50wsmwyHe7cdu0jhkj8CfEuKi5wtMnie2+n0
K9RXQrbf0dew/FGfduMblsyrljHQVv53VCj1U7OPoIXF42JWdDBG2dCMghggapPk
PA5/POxNot+yNBkRJHHi0yND1Okawi6hTQWGtmcLzjp3TaSCNb52kz1aOwfouti6
Zy5PifRRiZ9Fk8hEkwvFGhgUzYIDX+gLXcqa+gpcxNDqYLzWah6nSu8tO4/k6g7H
pArUt373/ryqjUZT5JoXQ6jsubfJekCybnWS+np1y83oRpDUmr0llk5mtjNwGJK7
ip1tVaF6Z/7dJ9wYK0axipB3PvtudYpW2k4L5yO4WUAt9GzTQWHv6Hul9QD79iFE
+GQZzaKbsTRutCaCpF1smGBE5PmHluniuZoyoWDHVhUpOODpx39gCpMrVCDLkAXI
02sNayyFuTc7Cb/fC+Xf03LHIKkjXIfvhGqrzHZiG+LA8wXrfMeRmEM7dK+f6hIk
q9RylBNEVB+lJM4I/SmiO1kt2L9yf10dzb2FspvRqbgVJP5h5aJrZy7qOMzrl6Ns
GzijlAl7cnS/IlM5rlTylaCr3TFAHRU9A6hX8RkYPNtM+fbjZruYKrrYTCheSI0P
dqlRKhgh2gnDUoeGeGWTdwbkU9wWZgzI0KovQMeffKAD//IssrxRk3D9agDBtnrd
Xw95VKQw1YQq8+H+NclmmZa/uX96m0oWLCECcOITRPzNrEEIwnRT/Pr0OdLN/WIQ
XVHzABfPutVDv2uAPxKoAuCcdsRR/qYK461lSDxRTClXB21Ks8B2AywpFH5MvzVc
JGmQO9UCi9G1iHGtJQrsr00I/PfL7DzJlxD1lPaasHjQbj9Pm+pLOOHibihK/VbU
ZnyMRd5SZ2rOTmQxljqS6p0Lztbz79hVTtoig+aRXZnnq9nMRi10maj+Ja6e/+Xt
7LBDDpzXNeXX4tgk+gx/lpf8Q4acToPmmBPiCv8F+mNQoIwV4EBsg+oSM5M0cVxI
bF6TQLppNtO7Otbn5gg+oKJ9jNK5Id8ENc5zT/Yim4c7ztbdQYDmWtyRM/Sqa3Mt
MbyIdT75UB60kzrifirGZoHD3+PWaoZg9g/nrmLmL9s0s/nKLPTh10faAWhlRJua
yxSpxioOdHVVZxS1ba4y8AD1yKyz1ClCsARsddEFoGUqETDmb6qLt+v/452GS5sz
MbcB0vL2wH0OpMv1S7rBWdTEeOQqiGoP31WfJh3EPy7wUks7WedOsjjfZoZknwgZ
MwDopltkrk/6B2NuWfKwu24j7qMEkVp0yVCr+BZxpY2frPS/j/zFIOfVfYdFyXU+
1K9wIqXV40oQBY6BZp1T7GMzwegRgzmSO/1C2BqKpVeyMQbr1Ao+4YieZ9/+xpk3
1v1tEI0eQwz4silYhfkuLbTcWL4+/7jNV9Ft6340vFpeQ64ZrVv+7IWuWeup+1Mi
TA/XvDk6iW96tXDibOs3VicLgQGkS7SfOscOpXy2C6n/h2jCEAFkLqDQqa6tGA9o
q9Zh1A1qGtoB/+aCdQ/m1hOSrFPRLW7S5FO8b9+DFgEzn+JWnNP/AZ7HA5ro5Y5m
MQPllwThsE9BIyBzS2f0tI+mJXsiUgQrlAVf2deHKuRAhwSGxJHM6i93fIf8WV18
wIS+pWv52NYRe9Ke0f9erAnADw7dt7decI7oJIUbEfHsbaQzLKclz5CSjOOBXro2
70gdUR3qFAEiot2+/t+z21mT8jmhtH7AO7Cjmt6+QoauD/Wn4AfMKMroMQjJ+jIZ
5u7WfInC0rY5cSflaZ0dVaOl38fVYt6W6adOhgm47JRVVFXyxOVAnTjhgzMy/x0Z
tPOqUFmDWMWvUyCL25d+YJ3VtNt99jNZRuQHIy0y1Rgw9REIFaoTjEdH7XQeDTOb
g/0ZvnBQ/tOPDMtztn6q6NuQbLPplvouNIaKFMYFzBa/wDF29WA0rDDN7S+qcImD
4yWtJVnOFYsLmERvHYVIuBNNEXKyrXod26ZjXHS26giNbTtaVg14sBrtT+3IrQfK
8r77UwLmkv7rQjQSj0DYpDdql/3f+VXBNhKw9Cs23QfgNkQCWxo40CmYFJsVUw90
VInArZ2lNIWiSfiDqxqWXJIYRk6vPx4h7n8aQhGM9rcHBWU8FCdgwhS47XfBBron
IzHZj0JwH2rL/bS3LYHuG8IXi115fDX1K/4glfFE8+VJNl59gCW2oWwy4Ttk1dQ2
I6NTMLL405ThST7l8Wy+tLrMzzRfPR3MA0yalMmixuMPGZO+4ncMG5UwPzoAFTlW
Fvr50o90rebz6hJppgaNWuzYNqcJLWRU4MmFgscL8fzm6pzPUdrCw8Othpr6pZmI
d09jFVn3zDClwb09iH6iqQHJxcqjldsdanQPVKnKJQOFMwb3fBxPPOWvslA4PCuJ
dwsWe8N2U0vafQGt23Kc3WqJEzCCym5NNRcIrFRwp0Me/CahtUz7YWtGBXgjAwEB
2LRzSTlMP2UxEJ04swkFO3cEFGGEr/tEG5iC6JeHE5VK8wpsWZLMuxzlpbWRUc8S
Wpl7R936D0+xaKhaEdk+tan1BbsdoQjIDlHqcW9zOGw44nUvfnh3X1AX8CQ8SGRY
KyGEW6UYlRMWqrqpHhEmclA/Q7mnXbKNivqqQH/360+6mrNfGdXqHG3ma5eBpxHE
TLqWSkqteWw9s9885onTPD/JHIps9zhjGnptqOEaztKI6QOwPXUqmV7OomlIkPmi
WLejdvdH44pw8OquFO1vrlf3iZDgs2h+7qCWXr6CXv3H1iWtzaieI1W2tRDirK/H
L8mJwiUgIPS/04sbQC9Vog1HQ3rRezTV+37HQ1cBKwtdw2JdNhL74PrGHINikhQY
qzucJ/sQMSCA2dYvWyDiP0CFFvtHpFUFJY86g7qcseLlK+WYoIGxyuAJw0OQJrre
kCXSK3oewXzb25xutm7uap21pScHs2wdgV81Td1LRc2GygAsgvrPUpAAPxrJ4zod
CiaFBga9ITflCnzr35EYd5CSReymBkIh4IrFLztfdqWyRr7koc5ybCtgcrfZTbxA
nI33imeo+uLGGQ6mos6eWvX9t9m+COwnZTSQ8GH+DgCdnrqXIm0nX9TZMcTG+L3b
zX7Yg60ujd1L1L++YBrwaMg1kTydtzPvvfrFQFY69xpHGWg6HoJN7nX2Ir7KPIL6
XSNO+A3ViYm4VMNYYjj+Zp44eXnsrHF+Ou0jvxmMY5iuuWX1WVwygrRGu/DN8zjT
OHPUwYftwAchcHctZSK02kQ2MUIHEZ6n3CkKbwFifoHV091v4RNN/0zZFws6rGXM
yOtPnM8+Mp5x4gA/r0Jvl3qg9H5cnvWP6jjwdsBiSryEkwVV4B+3h6hxkOAyHWeG
Mp11UkrOvhzJu6WS/KcZHnazOvKtiJwaBu3M9OHNJGcRBnJvMzdpsXqOo1IHxx22
YkklGCuOaV/UncLJpUHSBoNNCCK7XU5x+//V7SuajOH7Gf/w1sU5Naoa1BDplHcb
h/+xt2LItOZIr5ypNICcjwvPvIGpq0aKib3V9ppEDRM3KxN+Gy3ArDJ7AtkO3N1G
re6QAgzFjlVSpJLPoF2IqwvegBnDE8Vr8NiBwgP+4o8G22/EOeKoEiTkoTU0XCM2
E27M4T/EI2P4BKUfKZOglTI/zZDI8bBQsErm3yCQMOTO7xLe0ACbVW4ZeJo3ssmM
/p/xYOgBdJyE8s0SRGniS2rs3jxbe2+7cspy4xg0f5/UPtN4D7b4DwU2CWDIDm2d
lTqTclG1bUGxkknYcrXVlA/9ZVzmrHeyaluqiXRmgaRdSh0G8WVe6+4GATIS+aXx
mqeoHEnESBf56cO4r7kFDYKOTKJKND2hQNAwZx40MGhpzM0yfDPz1lYykMSga6l0
i6TIMVDMFD5sGc6hvGqQL3dmb17NkhrFF82DryBzp3irK4WrCTp4q8aqWR0+meus
RTkGnK6qmDML0g11c/TRKiSMCF+J0CrtnFPMmdNPSs83F3GVarutzqfYY8icypOF
U8PFZpIPIBBC/QSKEzsXOHgib05BtAHr0K3o+31XsLYrPQWdE4qSw6X+1QcDH1QI
WLBWc0MJwRhB+Go73cV6kCcGbUs1nq48Qq1obSpny+ZDLcxBYKJtGmMh19Ixaiki
9XIJNIcEH++uR4aVb2odJWKs9jHuUw5lc6RdIiXRU2xf9zfMTB/fhYw/ueGJoBxf
KdwKOlNgVQfMP7HNjqOGQVJUCwsp9zkuDmaY9sZHK2KwmCyVIE6Xus3KKZ5xHG8J
tflx/DkTZ5DL6TeJMJx0Lxy6U+uWtLfh88hrkj6+sw9URx5RGNPpooINOJzuz63L
86v7a3osl0q69aU//ewYf4mxc7pqPnXHwzuDMLVfWcQoHeIc47zgkTLXf6Y11a64
6GBx4Dvh8InUMRvo6BC9BjBKcj0p0lH5KFv8MLOUYRGL3i3esOQ0DYVN1P3o4gK9
pDhf+XhiaiUequ0cerLOzokeLh1rRNPZySGj/7jeN20tKrxgpSM5Ot+Ec8C67qfV
X8HlLm4VjXSYxxZDGc+mv8eSnBS619lgguKDiQum2TIzZXLKanZIJgtmTWPA1Rk3
IXS9bL8qLHSGMnS1JzTbdFrgMsuKbgGGFlCVomkIhQmVBCJ+EU7LP/VD6ExdJUBa
TSqwFuNJYGFmEXaRbMOePj041N22iTYKtm6lUjWrB0mdR35HPVGKZjfk6PipYB3Z
EgHneLlBM3SszKkGW12yX+Ti8+uWB5TOYYASS103zSIkYb7KCqGrsUDWjY6IaSHe
DkMyzSh6+RmNR5IWYCR7V4mAXyF8S6ZuUvckZjcQzr9IMBUnGUFL0EH1ILe1G8wx
MMuENki0XI8oQ5TtTkrtMxtaHBbxOBQ6NYeqEy55eTl88TqLMRvj6PGvjcuGITsm
aklHBwzFbPL54x899GZPsiJPdgp5eyG1DVAMfZmJjW0gWMHybdaj7XNQaP0qPRdh
ldOsfc1/0BM3X1lWUT0tpo7lV7X37tgMUBZ+6FigOHy/4LNJtfIM5abWcVaEF/rl
oiTUK3gHujz9v9z3EWDGhx2e9QVI03TVcUwRM3jI1OdZQS6f7SMjSRRCeAgndUzy
QaXo+VrZQ0Lm0I7E7pHcnGpqH+oVhSccXlg+76+OJRyfB5wZbUtFqB5UjT3BoqYH
`protect end_protected