`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 35344 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
YachDS4bpHRDzLXFQC4CtegLaKNOhJH6RzXDGQEpFlk5nEj0eTmsWTacTi4u4Wsu
gD6xil7S4/W0dxEI+qc8g5ZKxTYIR804ShhwpoVFWi2ZFz8yUAd9BuiNpugjG1oR
G0hlC8bzaDwUwyo7T1pIF+n9KjBj5ECe4viuPokKQDF12h2siALyz9RerICuSHPU
0Bu6m0EuGRR+lo+6YSbZPSDGnZdEqKnZg2cS9Sxonb2g5Qgw0r/ZiVGXFwegmAFM
kbzGaVhn1W2ryZfuGXVhlAFP7uz3sQ9JuY4yNRZ2HBKxkmKU/ptJrUsZzrPhD6Eu
mhvhtMCPLM+c8V6QD5eAoqyjZ141xh+WCknmmBUkPGqG/8alCw5NhMJdkAwKLAlw
oYR1gM09uoKGb5fjFZpzGwC8M8ZhJJm0qlMK2YMqWUPNcOOeAHs0LTtM0Z2DPwBz
UhOMDHGYDh4/Gi/+cfMVtGPPs5kTf2eAstFI4Hvsj0tPXa/qwP2s1bI20/+zyOKp
Vmgps6lXWvCehRfvxmnIasCc78vqiWH2LCizMtLh+a0EXhhI9PS+aRbfuY4wgQpX
OBS3ktr9AafLrC9hB7d462c4YymF62sMMLTXsXw+lIR/fF2G1IbzVaC2s3YNa72e
sN1xTMRYN3tY4hwn5T4rdszZ/b6Wnsm9Lx2eGLpFxTbIGmYPYF7pokSBLozmdQM9
Pvy5RIbTu7VGy0TfQflK4e1VQM5i/Za0LTt+a74BBOMGKYmHqBg+J0rr36PeLb2f
Jo9z6eDdDhHOjI9Dy2ggSXwCzNvyiCZUcoWeEZTzD51/le9iH/B3OAl4t/m1AJUX
NrdPo/PjxZbneJn4KQhQRp6KSBXtO+EYdu5nrsbpvxV3ZCcGXcOjJuonIf/dBkqn
BBL95ncteLSxApa/uC4oZa9ED82R8tlkkwObck4x1/1R3IjXNPQdqPgTARBVyqJU
OOSzJDZHRVN4eWxNczekWW4TvGLZAajeaBXvJiy5TZmMXcQZOoRatq1W7YmJqkJp
AI7e+QxXGVkG41wxbL58ts9xkSibjqZleoOL4KI6UG+Kx75wFO0Qog/VHSQG70Y8
8bx1V2mjl5ehzFdVcjK5vHPv3lPkrQooBb0qOtaSe+ZKJk7WNrh19lqjJLHUVsXz
ucN/B2ILH8HS2NKlu1sS3tlBG4+XXuwRltnimeNYJBmS+W7EMRdEU9Bmd1g1fQu3
7MO3Tk/8xpBMJgKyBsZ7lcPcvFVDi05cFjom9f23cIOKEVj1XbASY/4YZw4U1/fd
v4sHx5kKchj0QxaEIRzbEyDOGGzv3NihcM3GxM/ryXTcOqWakE2WjsbqJ7PxItj8
tMuZoIX+hjoYLoqLdYIiy4upJ+MNJXLt4XJ0bPp1YeV4aFfafFikmnEaaBTUmevO
9ArOQElD4Tbm5z+NMrrV9HxLZm7sBnF1cB/uGcQzUaRbt+IbP9uETItjm5SkdjG2
5TWVkW0JTRC2AWVyoKBY1CEqnBFIhslYwe0u7O4Dp8n3tqrcdt26rvmbD2fuZCrX
E5ST+D1tqj6KVMdj8tn3AqLCw2jbbYBBw0gDfimHYYTmF8Yo5SjEvb5tXUknVlkf
VHTjrFy0hF+be71mVSMxNJ98d94KAD3FtSCdDAVsDpymeClx7txqhlagE7/5HNQX
dz/psEM97+P7FBONgV3zMFKBay7HCIjCUIM5Hp8ugaDGGCFkc4t/t8tkRpyq7qpV
y9HB7YsvEYGPrVCO57mS64/ubbFLXWhF5WKCTX7jFIqLLP1YAaNkArZXqzYGF+kd
Wa+z+g+XGh5L3J07ujWmAESXWHi6mq43Iy3MyD+quSXiisu4kVNr/gGkNhtnGAtM
SkDZAMvL10C+W3wRmsNl25ivKcKn3mNOOkSIoxAfehcnuymy+BdTu30uTKw6EWSg
6UTRSrQ1V56yvfLaUM0b5zG6HTrr1BG3WetnRx2TvDa1Wn7BVePmcsgI7fYEsBM8
YT3l/aLWGGdebDEXjjUfldOr3M0BrssdiT9vovzVaaM+XOPvtMyj/2t6TN5YYrLc
a6l5Tn64tK6pyvSyOAVqdmNe1YN3eDWT3lHRBwIT47nEuW9NaBbr7rfXIIcZT9ql
sRy+t92lSbp6SDATe2mY7mR4Ajg69BkqzhF2XF+sHbClhS8aEz0WjaDa6r/MtLJL
KwV+eejUyi6OEjDY1qLBZuyN8fOZXLhC0o18GpKqVCMq6KvkJutWH4RT2Tare1U9
mNEfv5elVv6v7rZE53FAcA+NbaLgE3CwtegW4ye4RCRlLQXD2MNfDcRolMXdzgFu
19zJpMQ4x5NrhScscoPNHwAK3FS7EjRUgp9vZtXUzJuX2d0MjjquHitlvTRmFyMK
R+3YVCWI+cKNL+ClciWZWK0vBQjI/CmaBbNBiTSmmTgYULNcX48uV+ZcnUA/NXUp
4x9+3qKh/vfr8XhSr1D5PfLMgHUEMqSxKkJAY4pllVz91b3rnYoVdYaiqdyjmYtO
UOBT3DEHM0H2uhCwGvgnsG746/Ykm9Gir2VKPZRiKuwiEI6TP3sHBYT+BEZ7F0Ni
TqciIYCEyWR0nVYZHLN4asRUwzgPRe2MPCEc7A1kXtSWsldNZc+L8xVqpSpUjhrJ
1iF+CLmA5T/3ktCwp8mddBOSOyYeKmB8YhUxn1Gdm5UAxKKFG5LlKn9YpKs9ku5d
Gkn0GpfN/zTVdZPjq+leYd0nWnuBRYnZ3l+++rggZ3iAmT84IoU5LbtR3wSxoijI
/cQzVLjYhlxt8ItVwUoASIOSOK6KZic4TYNJzj1qAbxS7J5Bsld4JRb0sZj1h3mv
BYUcdWK5QCowyfHOAmPMN7u/jplKt3g7hxE4J1vvMJ9rYDdhms7jraDLxQZHvleu
YSOJX1ZW5rU0GehcH5ueLocz0ndeo72yoDd1nvPRtBo/8JqJvnb2w2lqakjAgx7E
4T32UujR96/lPXYh+coEiBZvSf90rt+biHlazll1WaTzHfq6MxphVEFFa6hH53TX
5iq90KWTqSQMwCitKhep4Gq2514jR7kFywMsZrVmWqW+AAHD+wT/2SI46KM+gaUY
8jj0LkyLX/s9jRMWjoyEE/U6niwy6AstXWynt9/lP5Z6w5Q3HXW7QM10pieZXy32
gUnPDbxmD8ZRXYKd3fqezXhM6uR+DfJ7sOUI52Nvqbdxq65UU6LcWKnTnCBVwnDb
C5lT3SKM7U7/g9dd08GOhNvZY4m8yh1GFWK+ARU1QqDCAvx/yY/Uc4+POx6tJZZn
RhQzhgytM12cJECOiIbWtNbHNbpoBGNjlaOJtk8Dn3dSIYrtEkuVW+GQNfyae8pA
0yxshtMQsFSgV5kkCmncWAsByi8Ozq17nuPpbzkgvGaE9yvFrXvAMM+5Ecv0cB+y
ZvsxFqgmU/IZlr2SBVgL3e4LIjN0aEBUK+8O3l+e7uicG0qJX6YCNGfsznT8ItN3
XGMCn0M7g24f93LggFoWJBd2gWJdD2N1G+W2sGJAtV6Kuti5PfQ9UDscruzoMaBV
QKxpUrHoqmSNLrk1oL9RaQp0ZprrXIyMJ1fj+8JN3prtoWC5g0ib6oS15OllTiEw
FvmHpogXggfcRfYi++eaF448Xyf4MsCar5VT4OBKEpsgOgfFaqgPhEUzjy9yQAA6
2jOsvXhabpkYAt5OXYj8peUgvCE4Vujj0u+9EXEX5CYjyI713ICNCjpsIPna5tgS
ofZ1WGnZ7nOU220UnmIQ+Z79+iHkslqVqgPdnYKmG5bDUc883LGNRLLFOMk51Bt8
LO6ZQJMp0G/rBrOTA+7mbW98FhIHHd916wdWxq4e/gag8Kuu3B2sP4p3TIDJEKVV
mwb4loh3s0Ncab0znOf2aGwYlgU9DvGaMAqKYyVFIL54C3h1CWM/xOTO+2KMVKSq
Pwf9NtXG0/vTw77VIv3brYjPIuAYMV+cbh42E9qdtDzUYmAqvwVrqH8Dc4V5cD1D
43Qd/dt2dqksqC6z/UH7ahtN1xMVCsle4yfyMyNYKL2/Xa38Wv35Bl8dl5Pf/UqV
gRXhRtMYt3AQP9+Bh0LjktDTlb443OZcQEvCLloqDz0WA+joIHyKaN/VNOAaXLS8
KvctHiVhsWEAFGZNmCMwin8slbSfz3gI1rI5oYQcFdbGmX6Lp1nqRBTyxrXfcuGM
Sz6Y2TLUjf0mOjLxjtCmhFCk9bAiL6AwoAHiesJikIrCJPml7dlvGa99BGVSVaGU
3U4lteWvp7RM8/TB4XpSuOyQd53I2oTGoTR+cXgdKOPWEDRbDo33Lb0/Z8kuk1PH
UdeZ7lB/z7v9YZfaOjgyfmyFKz+85HYDhZRCerYWst2b/RVt+vYTYQSjtVQKECV+
umMaJHGtFGwcU1JfMa8Zw48xnAEqDUyvoIEDtWNswgOynzmKYa7BQ6Fiadd0bRCT
8JMXjcfAFpS6F7KZhoTQiMFTQp72DNNB269IoUdxX+T0Ze+N2wV8U+lGpR1HtUdo
vyox/CMEepc16mED8VP7ojN8Brb9BmGKHSbaNTo8DbcwrWTwovCucHwYGbAxh2T3
P7bStVx6LgK90LrF8ecOu0Fb6az1jv0lXkv8q+FRrXSHeFH5dB24PKaNy9D5RoCW
auw89tRBM4JvLWSJ56op2aFH0hI/+rbVMMcwjqx9BHFOLmcF66R/f0G/seg2Z1aS
vYiNfx0vOKaGj/Bam3a0Nkjgn+qtBPtAYQoGhxja5YFHBh+MQqy/kZHvd/iGsVr5
+A56gm1CZS5dy2Cr1hZo1VDL5XPV2lvp0z3ThdnR+64hbF4hnwDUkceskujOI4zy
pvTyOGvCxe41qFMzaLwDR4ZcNcif8cva938UuUo+rUZX9WXKVT6dfaPbPWDMwJdv
9nLKfrumjmscI1GUcLmOQwkyhAannTkbWCZ8pQyAmxAxNinmQwn5HKdiDhsTAsme
bp3mlHU/OzzzD+ecqaDXRDh8H77AV3DUYPwrEXgPbmS72VHI1z46QjSu6gJ+7sQC
jFhbM5NjpWziIEBKmr7oY2UzhrNlPYpSEM2KogS/smTuJ9jFoBARbilR92FplNJk
I+K0ffuRVtgD0/FzSyQTJCgrgJUcupcqfbVr5jNuUu1/41F61UyU3OGdFuxJw0Fg
PAt3E+C+io0fTSixdB3KkVirjF36wBdlIHoogpVMNXDDGXSYoxavso1fCfW6C5+B
O4ioinANuISdXF3uyBCo0diPZSjTuXGqxZQDHb1/cQV3O/WdbjvWRF8W8n4s/wIB
3U8H1c+ELgBOgZIA58z5RCd1baoOLLGy9azWnwTh3bzgxBrUcpUKnNFw7JaS0Vev
ECE6GnzYMCVUy7XJShHsFMcnEhisWtVQYzy4LDXO1zQSqYOViwvXvIWg4GeclR74
qdNASUETyNuqCcY22iOG/UkISbBVmWdcTd4L+RpCvKtRYG4J9Bjm1R3I+ye2vaOb
cj0mhAWSUd6ZRkFZw7ThlFeSi3I0vk2cun0S+4fYqtHS9A5Jf62SdWDZXiCHJ3DW
gIUA1VK5byiXFZzv8b+3BmWhxQ8JE28eXqXqiuPQJ1JBgbuJ3zDmBWMhU9y0j+qB
nT68Ry1XuRZvtKvh7Z+qMgrYqBSvJnaLHP+eDRNdUL1sktZCoDOy9RaoAuyaiVsJ
jR8+FHPknIdtGX/68pQPfm2XvYrDA6yWkCOdy8qgkcjfu9+QOfBpxE5/Eb0f1Cmv
8ZjPjrhiHAK2n/1jS55dUl/M/xHh7YrqonlKhK2rZh1ODcvEXRBwJJeSnVNXCnSF
hIJI28gACfGg92OOzPB/XM7nyTZEdS7h6sRWxgaHYBWg4S84TbWE6ytjQ7IuZIgr
cY4IQVNRq9LhFiWzvRAUCejRHA5pFLQnj5qqz0VkcdTnIjKslXau3ihY6Kk1OoBO
SnNsCPfd88tmjkOwV3VCXhZi5Y3SRGPQ5PSChMIWiDOd6pRLDdo/uclXWhKLVtgp
KMZNA3cXIgFJDt9O96T6nPzNVSMUOrUt/6WHOlvSpoaHAbmoA7/mhKvdsJn10Q3r
F5Q1UXtDZrZoRHhlcHRzXatgwbO02gGBaj+BEQAhrcp5VsyQASskx/5t4TF+7+TG
+Eha2u5DkKNCI/PFGSTvOIDHED3Ute+caWgAgdyX9ngaosqLJuFVKa896bWpcyiV
0YfvLa3VCQw5mwuZikS3b7OZYu4Ksp8kAyd30u50PmbOkYNzMiqwNX4KE0QE3CH3
crS83fVWRasq5t/aNrTzzY/UnaqcbOBGH8AIp8T1Kee7ZKZAFYGMU1IVoO1bdEsY
wEjF4lnnu/fQ9+BU8xY3IDmf0M7tXDRyrfDPDjDqoJjtIANsXLzdP0G6mHpbR9rU
OeTTV0T/w2YhQO+aor/bNz1as8CpX0PjSNqg/fG/7PrGY0qaBxFs+RjwiMHTpWW+
Ea+9dLaqpmwBEn5d4MLHY0RmkfaHHO0bDu5JdfoIfiZg8A4Srk/MfPGs48lUnIfQ
UCH0Xv6Hsr50AbuMOXe8NZ1sb37SMMAAjGBtLc0b/j7ienlioDcWI9E7ChYqT9xx
97IyDwINlPbT66iK28nPbRyvQH5fFfmkcFyFBHZcbyf0gGtUj0DNh0YjZdN+xKUH
qjnD1i4r+xsJbXLIdTEPoNfRHOvVI8ek3tNs1siJrDoWtJ/YIU3V284LZg+W4nhn
e4tQx+VyeyZcDe5+GijwQZ0Gvlk50ksgyjt6BLYVENRKkkd2l2HiIB/0Xzx54w9Q
BiFyVNCTUt2fjl/Ip9Y/2Rkw/V587Uj+rgX+hkHfMgf1yQomQK8C9SjsuHADggWC
mtbqUYJuWBhEReJvS5RBdfIqPXMieZTG8coRJCT6cPKV8sy8effUev7hwFYtTmGh
CSVVtqmd6R9dMdRClZA/3pwxAf6WCzMoazyq1M2eyv2N2ToMarXB3w7RfCq6WzKq
wOXr2QZNSdlfiKVKLQRsXP1p0OKy6TmtkwLxWKbvhR88mtGGFIF+2lLvmX/c5Mm8
NcKbOUBpj07wm7neu07nH5OXJpLfQd7lNuImoNOpwKrkeLCJyUu7WGLIXnGQWdI2
Y6QLoARMxOHwx69CaOVoM7++ndEhR7fW30yg6upWnAtse/NhennGs2Az/0rUHLq2
JsfaK69WwmQCis4V84eMBEMMNGEKbW1mnMA6lyi2HDTeiNnm6OzcrvL4zXfOvYgL
RJbJrO2VMoMJaB8/WCbEM1HQVeurMKdfg8B2EAznofKZ+RBwrUvbXTS9geiuaqyb
Wwa40u4TU5p5BCPNv+0kcwiXMF+dt8m+lC0uvH5euBKF4zfO96uiqYQpbUVlq2Qk
mM0axY1hQFhI1KrF1obh57Y4BOkAydF4X3yoI5rMX1Ympz+PZQhQ6lIw+H9CYaG5
uWzbqZyE6f7xxGj1wJ8iIAqR5HTlCNhvxXXNABm/Ge25N7JyRZ1Jc5wb8v0F8dUW
GSSkGbsRpO7+U7RQwubW2NtHyoxTInz9QISxCLBj5ueY3GfybDoMQzTflNIwmHMr
qAFFvWLmUC/5LEyCqbxpF5Ser/813YcJCtxAUXmxzh+rf6T6DiC5MHU9x1atlVLP
Dlymcch3/VKL+bz8pbU5Gn7v3fBPBMnoEGjMhDZG1uTjwwN/VLxbJFc0LmUw0zB1
iSqWoanXKo4GVQOQf3iQciDV8a0pZjMRsnWL+YcFqfbMcjyyr6uvsbSu844FDmx8
mPL6bxu2FHQZwc2WUXJCz1AETqtAvzeD1vBhvOMe1OyV8ejx47Z9oaugzc4FH+YM
Y+tbyi3f7C5Bm7I+6NQPLMFVkeqSK9HZPrWNppKJ/2WaJ2pytS2HOm3KS60vWTZz
VP295A91Oq1O2u5Rsm0MnXSJLOrKpuPyoZfpHFMDOK8hHAuYWHNl0sgpvlz9zbvb
Yo2trAUmYIXguqwt8Ya/JCJBVbk9YWGRUmgVwhXk93P/958pg255KZDUwCBSykQq
RQIkb41ncw4783+yNpjcLukD6keQVx6TxSWMEVmvMzgBylbJzqYrPX1/3Prwmpnt
VKfLu8ThhgXB/yu6xi2GOg8Idd57q0Rl6b6fEiSLxZ9432FrU2+4CrTFhqlmX4mF
6BaMAnAoNMUTMbyE+CNTkGiE4CtkzFNiBFvWi41HErtmGPq4uyvUCFFxUMMNwzSz
rt7daIIDub+tJ8x1G4dImiVNBCw/LZkmeeMoJ6HbxcRR0p1LxyROPbUib+ShYIyq
eSR9TJ+rNw5tkDyt2OqoSTzqATYf8kjGQW6fSEq6MddHfRfg8J88UyE0o1kRVMnx
m9hwSb1vjXGymZoTotE0TeoULxZM1/x0fxyyWUVJSPYW7syekgSovQQZse6G9At0
2U8fPqrp2HwcLNoLdqxUGAV7LiRIXUPm5ZhrbMkSf+rAqT9EcADzL8sKpkTs76ad
6+0lwxu12E8VVSyJCTnSelsh62DXFDV6eWuw5qPTg4r7UEBo5Mz8q3ErwkGJf4bH
TdG6ynF+bgv4a4AXJiFzzaHEXznRP9S9scopB4SL7Guvm09KMZzP0sO8p9NY60va
0HegIdaBP1MbDQFqZ3gwXiff+EupSdgZCm+5llBd8ZEdWkUZ8Rjmtxk0SdzrdKX8
ENewibm0JMqTjmoV5TewTwF9OspuYUum1Aymp7PJziDV9a4FoyG9FBdb+xSeozY3
8T62SAFOarJ3RPWXbFWwnIshmtR1LQ+w1nKnGuoe28feNOVvUHh2lWNqp49rGeMu
QiHXPsKuRufqQ5m9hCtpdzaKuUMOiGMHLRMHUwv08VufmN6vGVB4RMd+1E5IIeQl
ja8HgOBZl0rOCvLa+t2NcwtbuWWv+smBnpTDzcEjE+WyhFTVVj4AG5GbTwYPHqzv
sJTNpyYoBdcstHe7u2SuEmDvdoASLXushwttXlt/Zr4IQHZYek4GfjqBEOHipq7N
E2n6ACbH9k1dLbI3AOxkolYeVwZRB9a+yLeYMJ1lEVYt/Pg6gfIHUmeHVZ9G5d9V
yF+lunHoM4/9jCGkEfN/qmsvgxt6jJZMHP1cvNkpJqxYuJKFbEY0HYEV3dYAIJE6
hSY6fqHFJ0MCKC0uGPnrjrzOTSEkOzpfyPSAYyMjrLeZw9smKhe2mF/U0j9ogXCQ
AqDM0GbSLjacQGF22q2igzZmZc65ED0U/ragFYyOXUQJzuUmaP/8XhRBj7Zkngcu
zfOiCRj29IR2zAHbFZiubt7feGTjvv84e6U6MUkK3txZgYnM+OTXKFet08cx/DoC
IHFkw87gxXAklESnDiAKfZh/DE444G9JQY3C11eZ9mrR/QycInl0bj9EQb3pis21
yPviTHtWMloDOWkQzETNQcKD82NwOYS3BhvINVqc2vuGktJiKaAbAAUQkltyJ8d0
x8Mi0hE2A654Y4fPrw+GsTou0mxV/+Mn3qA6FVuQ81S6m9RTLC0mLmtfy3IKxoCt
gEVwaQM++7hKfObmK8HD6B6Gjvrce/vX4JieArKfjDhw+pS/8S4oaJy9LqW+kD1l
bS0XrGvRDB88yZYlBDHtPG12XYBZEZshYN3uOq26lo3GA/z0B5x81ggUNKbS+n6P
8IaZLOM3GLbiNugrL6TvMClereons/i6un48rEJzDtjndR4KXPWlDG8vD6QCfYHr
rUmqdqmwod/TJFUX8sOajXczl3Fyto0VcZR8KcKqTFHtaL3WWLsDNs2KjMx9j3NJ
f5L0AntRDbottOJEIAx+Kw0snE/4Hu1lLxOjo4vea4FFF6S3RtNLyEbzSki3L75v
ZAqZYp5krilyfI9VnaPmC0pREMD/f/1P0pM0w9bILXu1Tja/1LwEH236qtvK4DjX
/l9I/uZeTfahl+YfQiGy7xqaNqvbWl55MLLXxOwp0DQ+x710ZvSJ15ZOSUsvF468
TJqzyLjqe1sGFRlDHURO5QNA6QCKcXOZs73mg/HY79MWMlrOu9rFTXgC4xkM33c8
iSHnq16+7m4kAsvxlqM28oDvNOquylXtRKvQgyi9MyOR4YqSYmlcpdoap2IBh8Ln
tJ5UP2wHtSHeWlTzlKc5zgNpf2HMGxHP9K1j4JHXCz07lu3YuLF/s8DPxY2lEkCm
JfkUFKvhZ74Gbeod2UrQS8NsEYV8OxX4UECoWcs3wKGztRPXVSz9I9qA3C0ngxuK
GSNTz8dkCvBi9UGbQCG9s71c2irRvHJvhW2BPf/H55j4ZpcGpNYzjry7S56K278K
fCppOeGRTjpBV2GF117SmMBJgk3KgeU13fhytLdW7DydBcTZ/qNgVFJOugfxQBIm
HemjHX5qjVuiA4lFfBGu186lnx6fTzalFDbeWTj6SYzPuN6q6oBV1wpPtzxHwrMu
AQWs9xFIzpN+M+FJNTzgIPjDZ1HpM0/P/LUnjE/LI/T8TV28Syk/qF5YQkYr5THH
E4dx2WuAVdkaN2i3Ux85rNzbFnYCXmpKSyiLNBlNEIBW3lSA0tm0876C41pRpm5h
pKJYypxxBJuavpZmHZkneCCjRJtXnbWJLszJN/kAiWZ0N0O9gfYaFfOcibDZWMgv
ubsOhRMEX0vpxIFuUCZUAUbJU6NXP4nniEzzxjGyPYRV2h6RKKie7wEIKUE51Ucf
//y3NYbVRO/Ru5sK5I3Ky3brYHrLnkv3Nq7L7WzGbYNSmtkK0cOftshB/+r1HHgQ
LsnHCSoSm8hfG7+FQHi+leEnt/cEHKc1L2TN0AKDAjeYK+rvUQkMBRvj13KQ1dHQ
LPxCu9/Alw79P0DR3HGRYKh/XqmoeZS011Uu8dZjY6gib2eSswjU+ejzzwGEm4GK
6L0FIgGNy44nQQhid2pKXGGJf+b+ueqwmnUZ5PKzS1xk9dik315CxbPKKMvUPYZ6
CmXF7oCKtTr49teQTutiUtZT6DpuRNQQEtOo0Py5uSjO8rsbr6REY0aPj/XM5KGE
qeQPoY4nUP6NKT0asi/Z1XSGsy8UFhIGn+zSmTewfh0lK0MsIJFEd7au/RjnYHfZ
SmK/kq3yTSfC1s9vzSgIAJw161EuWFqA6insXdgaZiu3gLCNsJX/YAUl6lL9ll+0
VFlpo4XLQUY2CZnmS8Jh062lUmpYMPqC/HOGjUrEO+oKdMp9lTF6yvD7DePlKeCb
lJvKzbXxooGYnnZMKejnFupBIrbXJA/IQ+EyYLq0NMo7mX3nes1XRVQA7I0uPpeQ
jWftk60R/bGsdmnj58fFSGMCYO4XDWgeYsEcLoc5Oxigt8fXwcNnoMF7A/dWaiJX
SRYegg8J+Shcys16ZCjGqfXBG3jW/4OuuntLIIC9CSWbj22blcSo+WueDqvHJCmt
OnY24ta2TkJbTdA/7kukKDvMDad/KHsfNsztbMl0zgvi+LNh61B3YK9srtDhNUYn
PJ9R2ufxSJof39bD6eDwoVT827pKTWTRHSf6nMHhI2rl4Fdhae66i8clO/cNOnzc
5bQzT1yBMdIcgdgREr+nCZZvu+PzAs2fS0sqs/l3+4byVSpp8Y6eGy4TkZfp3Zkq
hgT4fj0IFBa6b0U/k+kpXyZ79LZ/VI9AkQ/O5c8mYmOy1u8jkFgyIDxwHnunyndB
WgttEjZvoJcFvUj8dyRuJ0eDgCY9MbMOe/WLWGTmttauW5Y52CY2RJM7K3mXeS6C
3CqYW2RBm5Q1J94P34Hb2uwcg3TWmEhW6W8c4eZfflWR0+rdb1K4f3VsY3I964+r
bYm1vyf9TuDN6QSjb6aGNmwahOyidiMIsyjHMep5H97sfeSAChNjt3M8ZT/vFsMn
6AcrX8rwLvFwLOA/61nRfWunuHqLprELEfxlI0oEgWiQZmxiKMFNXMvBBczhPZLI
W4XXvTABT/jdg0NWVZSP9BWZzI+vaxyhKS5E9EBYpiut4qmG6+rIS4qlum54ldRw
aKVo6FQnEMpROT5gQGhzbt1jUdGYkOWFfXqO04v+FlERNaYSWN6w7PsQa+n0f3y2
ng6awu4LCpJBzKwls7025T01mXDm1XDY5lQ3ONCmtOxUQw0ct9R+UO1sSmBJONUU
rJCyLsy2M8ROTAeblrWtFA1p8s7V3PvClXgtuqSOfxkz4HZrm/QBXvz+pTaKRkrg
dx3rO27jixceRPB0m1vks+Z7E8angxQkHjSM6XQmbSm7n0jKSkZdmgENetOMDx1J
ylAGDdvfZu0uaTBMgkE308BrgQ/8pn4Qu/FGmZnbL+1NQGkEtMSXrpjibadvFzfz
RwdxB0h6bcMIMW8ow4WIMoCYb/QZ4uaHuU3UibpRdgKTutAOAia83CxN3xeLCNtL
B3pijtutNQWxnB2WfsAzG7HC9+lkv7CqTYuXDAa6EqKOIFAZ5k8KEJ1FeCAXQ2p4
cPbVeeGWdthR+eiUBQgTyJfsTHFluESEra2CjshxtL7U+YpzTYHGZziDqwo0Tj3E
cc0iQppk/vRVQYuypYUCmy5yl2UlV27AZtkPFzML8TgMmDsKCpoXsCJWFGcOCUhz
l63a7utrnw/r1EzbGI6bEz0xrUYdRfzS15DFUDwy+oEtEaA3GFPGnX64lQBrcdyx
wuZSTeaa48V4VyPAtcRS5eyxVAVy2UaQap9m7FNjhFv40q2twTgnzwSmNBu/D4Lh
9mDVQs6+YlZY68AHbXCRkS8O04DdBh5LZGYfOAvdoEifVpi82qgvsSGJukTMiMFP
Dulw/+9XKhTPSonp5zVsJIcb3Ylc+K4aCUeuI9H9GNwvcF+FLWP4fQQM2tuqnkAK
FnIcWed4nnXFIoLRlGBsPRN9zaWtgsV/6MH+tc6UiG9M/4xteE7syrvIPGd/zYET
2yUcTpr+PezFRvEDwGbqIyyrdQaK8iJ+KF6eDRNbE5QP+1upaijsl9P+mruwuti3
o9LQXtAE1GiXX1ZS2ydxPDLtcN8kTXUcJDgsj2g28J5pslceU5XAPd6RXSJeSpA6
rhA4DqADyV5xpFblNk3FnAYOnhQGxeTMoC5Pl2k7TSjGxRCA9g2OCKiK0iGiKP1m
q9zljKVKOaKqvuQuzWikU45afQRZFOc3QLkzi9X+oAgo6ykPbOlzMv8paRXIsb8V
XmFrIy6InrZEXaGSiNZYBarcz5Nr2Rp8jngfJQIpaop2tuYMLPJbAmxphQ0u/fFD
IrTxLCMGJDtCtChLW8393GMmiDZMj5tWL/GwrlzPRQQVtDU39hpQHoXNUCiV6LG6
nuqOLsZaospXKozKs0IG11xwDd2HShE5idDprsNRLF9+icnc9S+eQt8T5Lp+YMUC
maDElAn3GQRNjS9eACE3kUvdHzVH2pAzsPDAOJrHe2VIBVVQuz9on7vCkmU/G8CJ
zvNBumZomyq2ebxSw1t/Aj+oAlVoaPE0PO6ik0X0AjrcR5uQHtAYz20zvrOBGZwf
Lp0IhftfNrFlXSZRu/L42hGfDE965fQlitg/7Piwy7YEzk9uyp7Fqn43amgStGHA
0hGU5vg0FqCiLFhye6r3LiF4id71qkldWP+sJKe+O5kedhfjgIaDotuREH+Felgd
A7MMOOPYN3wcSxCj1WvMDv8ZnMHkTX1qMSHlk7EA/BGPYDV6aiXB025ILYy0iDVI
zyEY5vGNlrmeKxR8f5VtULiCwmNmUQcc+07J+7I2+ltQtnXydCTool8aNjUzdSmM
BuY0CHzRlhUVS8zqG6+riQTeyhvgGjX2oyp1thXVpW9xE0j4bZBoKct3d1j61xVX
oMzIA9TSEssw+YC4zLzNNh0UNM1cQOL4qTpMAOE8PZrfIN2mnhsfb1FymyR+pHmD
veiGnyuC8MC97iyneThdE1CZqDMlV8/tmVTuoSuqMmXTgsUU4/QvtUra6q2tV0T+
KNseLlVmRpLxq6lU4P+SE208zZPddzXvV4rFOe9BlMAOAlnHxNOmpSJASQKQR/Lb
hMHk+C2/Yp+aBICkFj50DeHGLrnA1Q5MS+EkWC0BxCQvMrYGgdBiyzT3TJeymj+s
ztRzErwJQm4no9hWRyrV5zFd04Aw1KDqI9/CJcMCFZOlIOFUGF1M/3IaF7RazT0n
1G0Mw2z/ljHEunzR0tI2XYMGPd+5vsaagQ7PiteY+zdC8o2JkPoM1dmwScCsU/gZ
PW0HwThAXEh8qvcrLUPg/55t3yyA31Mi54lGh/0YzfX4yusXTKV1A4KTiTIWRwxw
/Fb4gu2UB9zuLm9y68ba5EPfnHHshpoX2uxlUgr6hF/NbwoJYNWqXmQb4fT0naXj
38Z3CujJ1p+q3NjHGkzZnHu4Pgn/f7Pfld3ZwcqSzESe8E96EPNuibMVSaErayP8
z3q3YpoTVDG6z8fIat25bhCbFMs7qCYKKzU7z8N6KahO10n6F9HAbpsQhjM4TU1k
+HEy80RNReMd9C1TsXO9DOnv4vqP6S7oa4Nggx3NmGVwEtX9o33Fs3QHWGIzeR2p
CR4bA99FHgnvzNXzKtLhavKVpsxECvFDR2PT4WQxWYRrV50w6l+dIusIMHCA8cSg
JVO3E21pp+Xtjb7ab6VABg2MlOirlCZX30TDPStZffKTloXZRaXAbwHBtIdOl2d3
j8pO6AXoKUGgSv67VK+vwYNu/y1F3b+U2S09W99KImRG9BYUl6v+Dln4Ftmr407c
u67vOJ1CpFtUoi6hVeCzw7TZPnmkaNcHGiiRbEO4SMEgOw2C0anZgMFjNUwkiqr/
Vj/RSr6FaSs6NDZ60z4wpgLLXFwG483JIVisrdVZkv/z/mRS6lk4bHd3QbdcJEvt
/qHeCUhh9SRJLuEdKOvVoe2WHmsRw5x2LJ34+bN5z4ha5g/sV9z4BFioX2VBS7t7
85rawn7BP6EtKI3yNeGawfkv1CpMtSaJSMJWEUX6w6ZlsSdDgy96vzTxv8E8pJ9i
ExD1dtonxmhjMiAiXHPVNHpzz6iyif2sytylKdkp4BiHHCd5qYs/8qo2ebyVF2b4
o7lQw+fqHFVZQ1zPlPclLfIgj28dTZrzuC4JAyk+WYwLnJ8sNubBRzt3dTjRfZ9Y
ej3qGO6+9hvdMp7tR9UKeu1qWT5sbpaMZes1688Ai+jD+QgIUAas+u2GpX8AHnbQ
E3dL8b13Kz65pjzNQMZlP40og67YSdAIJFmQe+jImjECOpVFLWuf9SlxKP8nZR6T
OzwdwJrV+W+aRBF3WB+sUJ8e08noiL6iW1buPxaKJy/NCOZN3NvJYQ16cBhYgCCP
jROYKKqMTSRR8Iqdb5wkq5VKigjSXWnR2evIiBqPLr8lGW/4bhdCXR3ooI2nngNA
iqesFzCgP6A6NWf4bGzaKZ24qFR6IPg+D5yRT5XX4v06opoERhHkQJ08PJupvOuV
D2AsUeUgd9VauqwEKxklLIt5M5BetZTUl/BaDIhDssw41hxi+04UZrrrlcxx4Su3
0dOj7s4h045oissrhe818Q4sFuXW0hnLooyqycKkCSQa/g7xzD9zwgGYWDpRDrsm
vGIcuM1uFC7qfWz+XErrNj7AtaW5jTPRJayhKHSbvNJ7irS6AAkP1FF6DugxKHpN
yEnoaz3W80eeZmEUGIFK1nAj58Paw4yzP2j4n1JoZfd7XMEdNDUBcjwZRUGQ9Jue
poDra50DPQKLvHVCwxMdXcN/UBQQggx0fFgIVaiW+oS7LqDINr+CxqPtP2sAYCgU
EIW6aCBn2sQzBmZW2EkTeKTerGrMpKC7fynCnZtGZoGLhiQFkIPH2xL/ov6qlr7a
DhbPUBI1iRDnCYNTltlWFi/KS4wfzqDI7a6W9XgySjVmNusK5ZTJMPshy+/MvJqK
wf0N6s/vhhwKxG/IYhQN2hzEQD0uNyiHT4ceaPWkrtJsEJcJfzML+nCa2spIXyju
kt9A7K+cLdH7UbODTxgUEU5f4iZLoaInUlQe+tNTD1FOTM01NsZMzfmhw3Ul2gv2
r9WFrHNypnTJbdvSP5cT8tWAkDYIM/lJasKUW1RjGre1DLPi+4WVqLYoKtH7UX0e
MD1KjpYHwxV+L0bAqPCNRgjS56eyKC8h5rBP54drrmIbtQAoHZEM+ZauUS964g2E
AgjoQ7hs6QV4/FTPpFDf0d/KngsfEj6/aX/rH491WaVAfwmuYym376uWeGM+Qv7G
Wo5ejMfx7mDKyw3YnpGSg8N5y4yvnyY8SuHr6zQ2lA5gf9+XPHyDL2vl01Og2lBe
hwXv3ABhcMPPAPpDUnitgTm+8RrCjtGcw3aGswJxrBtT7LkP9Y1KwOrrPKVcbOff
9rhWaEKG9fM4LL7sqoEXM1RDAATZg26xhCSt1VkXHmvt80U8CGMmUvKdCGhCSSav
/bn7vBGIbjoCSY0nN/hSob02EEstOTlIjEK+BqFT7Mc63yMdvqamszQMIfzHC7qw
GZ5tZBxz8hbzQCzYSMGS0ikiwcGtoGZ0rw0fqbnttQM+Nj+gJaENoIT1apfAjX/x
NGsRjnYR0eErV4pPIC/66iavOA4pofr8yecQm+q7JH6LX/725wz+CR/itszqOAyJ
Dz6H4YXmvx58hzhdG0MM+LYhQntGDwBarCGvO1dH6ULnwGjIGEDueOHWvyiqzcEF
XJSvnf+B6vXuMpcXMDzuy2zNMVmJWOSb3Qihna/PY2Y+1ZaAl0E57c30s/b+NJsL
KX3UANG1XfwEE4TxHe1wZEpVOBS2mDpm7CCPOPhrkkyly/H5x28nh6s/tbJ7HMxr
gz0EALyPxYmc920yIeFQRum3rt5a45EWYGR3Fx81ey/T1sdifmc6mJuSJFpiLJT/
rTF905zG9u2xPEXw9RlPUeCZB214Jp+tuXji1HRQKnfHBVhehnBD1hpmq1WJ5s4U
gi9YfDd3z1BVNw7UHHuWmffVSI20LyvR82U3ay4vPqfDXIUVuPhLSyy4nP59B2Zo
dwhljLJoyu3m4TDwupLgrhrhq76Haue5FDrBXOeyf+/vO84+lx8Vzcbvy/qo2o3A
5iPd8iL/GtAbRQwIankbossXpjJjTckuebhorEPLAOjwqWAq0fX1P+P4K4aqhSer
poFZPYDJWwISjBagoGMSET7mb2U3NEk0WhqrXfwO+OlGy/d0zSM53h67qR8+ipAn
Yifk+RPa+L0e1BAw5I6IeikiD5/3l4/wWf500SnZcHaJG1z0qRR9eRr6myk7WiFR
22T2OpR8QU4qfv8wn71xALDNTNVgA/1/2Jitbb1A8JJjNMZOsrKSE1o+YH3pD2uE
Qa+d5g96v8M+kXPLelzEJBRAb4lr/KTIoBUaPZEQQN2FkMCwlKxYfTyTaeaU3GOx
n7cX8jBSrXXUnztUugqhqwjbJKYGZr7A4AiFk7mBuPV0LyE5cZGUW0dK7QXgaqr5
3oW7EzosxUJ5+p86HfCRvao9RCXeOhsWYME/fnMQ/PvQV9Y5mu3qNb2DeB+23e1O
kFUB8NClcqEY/lw/V1zwcpaxilVf9VSPk4/3Jw9GEYnroWH/j0ufbLHKIrmhrB2c
mUAvL1R+dbH1kcOk13wrOVuArsFCezGgp6QD6r24YXeMoRGrE93ToUR/IyEJ2PVP
v51PYtTjp6xILEQSeA7RiJh9K8NWs7cRjpdXb0kL/ChhknEnbps1B5+0ekNIHXbD
1yfXe+oXiYL0KsR9Q2FWG7nJ/oMOe+3cGTRZsFEtMz9QkkYSP/4SrLLEECYVidEg
sK1DEcJsYsT3Mm260EwSwwOzT+zCh6jVRuX/qj1KHTWBVU1hXyL34ArGWvY5DyCY
JVnPhutPzUXSqSwVVIRWUm0Hjeu97rRcIsAeJzEz2F+lc7LociHtSmOrawoopyXR
Yf80T5XawZZ2dPyOFVc6/lwqgYQbrw0/LVVw5zJqjp8LXF82CErmmlkjGG1i0U5J
hJ0KRBy3m9xLSoOLGUF46af3i5+XbxSkRAMwr/diq+2wMQE/if1NPXY9n0oQ9+cD
XjMvP0krRjoX2GLl6CcZXqjnjaoyqUuw+pWSCPRb0bCFR7g2ousqAZYYEsCxv32K
HNdFE+p3HwkxibrCcOvQH5j3fnp88Zj1aac1y2WkjdPnM3xt7uoIeB5TMP6u0MKr
QNErDGiZWgs7aV/Knd2L9rBUNG8CH62PhlgkwZ8VeymNWJqSRn/Q7D56n0g+4dY8
SWiptqQNCRYA7OtMaofUhXZLglrTYl2XZxs0i9A0GhrF8ipMjPW6pGL5/Pls3osk
WVU02jsYRgh7wjzE8m2AAI5NOkFv4a+3ty5ztwxDWQ0nSaft8wWk4xc1sDmY2l1Y
6+FACeZKUzzU8yBNHwz47M6kpDhv/gzm6WmmzI/Mv35+10BrtJhYQWm2AiPnRU+Y
6QyiIGiikxlvL+7fsFsv/d87HXqrOk2Orx1Ogo0GEAzPt5+B8xs6eo+o9BOx8PRD
oNV2gYiWeZbFN+lGngM6nC/G0pDUh5T8dPcIIlyxU/4imM03CuUjIBxPypp+cfjW
AMT0prGRhNuO3WJi/A6rOYLRO2gmmL2RS7yA9ekPxsuMo7W75JFDILG4CfuYrJzz
9lFTB0CbANeYNiXUl95aic4iA1tczDmNpwlFiqXPhSSlMDoWwxgHC33kD5LqRuuP
aU7+waLhnF4PT/6vxMpX6WFxk9R7SD4dqF8iO4XcQcnce/Sx2oWQ7j4bkTYfNrOn
xfAciu+8q4b9qUUiiP1pXgM6CD5AEXhYilThrqbd2P7ir7/PpKDVG0MUYYl6VGEB
zhXUWH8y9GYNRZPeoT3gj/3iWjVBf1hwafSuofouTgS2nlQcSvkwbqO20LtEIYuG
ymRdqbgblbynGslFcbOIGWsf2CWLxwZdokZlLvnEwHpD1nOIuLu53NNwzxZAKkc7
liF5q2wJbDO64qYzEEHTAj2we45SUvqf2lL3vKIqK05NeW2/Hzd8H8iejblRTuKg
Rxz3n4PoRLpH5lQ6XzEODPf/vdUStL6mRj6Bx/nraX5QSE0PcBKszoopYeqcixSl
L1/6lROK6RYD7s++mfihWVpWcp/QUWZsxAq2mGTjZhEwz4WP6ht+hUJnrHkaavWK
076jHg+yobY7DPiBA8ZcxDhyOFHdsJITomgahZatMF+aKHqfvRg+fvckMCFZ35uA
tBKEZRzp2qWUczhwvB0pFpANyhmrv5zCpdSZATgRwd+aLQppRw9Aqupf3yRCkKBz
TgwfJW5i2KKadt+bdA+sly04CW1VFpP9Oq9qHi0VAnAAOr0VCNr+4ctljNP2A/wg
6h5wqEgTYIbQq78h1SgS+AgVs80NW2ivrKsUD8YYXu0WN+nkwIO3digYIPySc64q
6+cK4hD1myvDlRL3UvwXX4h3laEfQ2dog1x3HXpnArN4hnZR18B8FciqdH9JYGPe
6gx3WZelwv7yQI0UiEMmS38NLxnqs+0xbVWP1tweUrEd8zI0bsj1gNfLwTZjYf2s
2Wq+hORP77q7AvsJ1kt9Z2n8RtEcuRrjsM4uRbxT5UsGobnclhjDYBqI88itlTdy
/5gYuK3fzQ/9V0pi3bYmQkWlPPH9ZRP1g5+KObBplLFuTeauIZbjFqyMe7F/M+Tt
PsYB5TUaX682JaRB0sfHiJTGVGfqHhcBxhvu3VxIpXou0wRpLRTv1zjB7qOXnkDr
o594Nz9WHW3INQyiNkD1cBgRSK9c8fX6klYS8na/9pdjgO9XzIsM/ogmFXkUfsKQ
SVe82vW6CPY9LV8/XHGC3ch7yQUtCZBX7YVvE+V8tEnkuL5z3KsKDpD/gTpmfQDM
YuaNkiDemwAjMlxzfI76zdbhx8z0UoARSLWK+IiXtgjRj4D00sDPrnE5677TrqW3
gbHQJdjEYYBQgS/5V5vZK3Daom5XhyEgPpZE7YR2oV0RUJB/dD661ZZeUDHKidxk
4nJDAmOPkc45mVdgpaJgBtQnylLXi9NWAXIdHfLdsucJMYCHm5mBFOf5jLC5ZkmZ
bvc1AVUBjETXfJ4pRpysjUEL8sEFmfX1HaubVaneN4nH4CIDdkBIv7wW9iY00fBK
NI0zkMeL0XgXTaP4XwjAeQgrTtWGnheElMftpAc2H5xuL9r+/LXlFd+HUdwsJWEm
L2vEvBbPAoOIMYE/J64zmECLKZ2GFK04MRJG2YUHzDM6YzxzPv9iRwj6MZiFItPg
yR0UU04V7IwUcTNZdTlLnJwE5YoJZf0vDQnhlhtiPCCwhRflYACce55kO7rISqTQ
MXBZ6R+uY0F2cy+nAZriQFJl0dl2/T3qXM/DdLY5Czc6F08J9iBhFYMb6ScW2YDm
JPYJ70FGnDdwN7otZJo//P/6YJxqbzWhXZgrr+QxPDNNtlcy1KuRLPj3V7pJBo2w
T/XpPhAnaASTq6yBnFZmWtiA8GNDEGYVPm9PPRPrXi207iG3SCNZBxKTZOPRF77O
NYuugs8Xnk1vjTN20lWFqo40lW5xG583DnfMu7LFp/WiMX7im+IDbAjsEGm1V5A7
lSsf4aNWLiL7p8jhiVElebRzbIa9r9GIrfseMvlW9TFbHFSyOlmT4YG86cl2qf2V
VFLjjWAgWNwzYhLprIb3J4awiCxwnumayBneqbmPgvyOLptvg6Ocojy7MtIev/rg
6+hQLxp71fdyci6mey8q4xw1JyJmvvz9jFIIKPjwyotdJ0LAQSm7aM6v2jKUmkpQ
lJuNad0RMknEQ9CfAjzdi0r5AXR0qMQpRNOKbthj491/MUSNSTKfbjMGLOY3NUPw
zKfCJpDN+yYr1G7AYo8TFffQQqqp/Ru+O4poi7w5Hgh9uvDPEhIUDIzYrmcqg9ce
oS26J2KLgjYtTkKW2/G2Gf6B+sgSJFi2YwDTziZJPSgLgubJlOVAtgjMRM1X0G8P
vKTlL211vqAsJ/jjWgp8nIGWDioBpePC4G68U0MIS4XdPyhofBVhxJCz5A6xTe1E
eAt2dHf/+rBvBL7RyjPN1iG41beqI0blCmwvjZwucEM7gUooTEWJDBwRZdls5owv
BCYi630VlM4CzWNjSJzeWodMye4wc44aShUUMM4tBfmjPCzXhQxD3UmH1uYtRIzl
7tKtwb27Rb7zlgXTjqZQF+cfQs6JWXmyNt/B2UVaEnBLHEHpDgNp2DJGTXZlMsbB
51L4JXSZUXgf5oQCb8t0up6vaGthihl8rgYvcsT2rXtfifSIuGZ1lV6jPbQFp38x
71feRUyuw3Xa9XXNOQf/wWdJbx1Cu7VVwxjNu64ufKnGa8n/4vEk7O5ag2Yo3r2N
8tZneYypQnm8eJW5Tzdhd7ppHBRH1b8Rqu7JMpqZ5Gk0eriLgamBT8yxbxP1PiBw
8EDOOnW0ia/IBWyijMGblsIVAg92rGoPVqbjBt7gIfSRmlzysSK0y6CW18Jp0bLC
rFo12T/l9Az592kDLGGaRHpeFHxrYqY/+CIzL2A/iXJDdkb1Odvohr8DCgSGuK5H
0dirwtjcq4phcBKGoFLtmSKrBqbFT7FZXv91p3qqJcBW5PkpdRt23MHH2HGEwqBf
Iw2wQNPRd8lg71fhRwfiH7o7CT9MGj77+R9mCqon3hYh79XoTSjUYIk3QZ4mVnhf
LAyKVkPHUr0OSKyB/10vzrmQah/ZYfxzbHLqnGCrlj2QGKY1TDc/xizsz1SKPjEQ
qYxpDKZNethE6ZVz18s51sAzWn9PQpTMm62wgKsxb1Fg725z6z8fqTa5nDAZ0Nu+
/hnJ6Wju39xgBAxHnPDqg9u4Yfw+u/ZcUmUyYeK82saRrgOV41TNbcb/O6ZMYyYO
k+H054x2JNOjDntBwOxGrMUp22Xo43HZNcM29drieQeOg45ItWfGlD97plivlmXL
HqV7i5tVeyacJbsTo2mCRsG0+mEKF+VSJmEerjK1OJw608xRTKeJ6N/UU2DnnWxb
+894+K5C5KQaVkgRinvSAVU1ZE8JGRHUgO/zkWw7KCQ7IKdgRScyB3Su9IQCGlq1
7jdmYKXtaswvYr/NuVf09/U3/TqbKT4XFU/hRh2Mb6K1nteuLEYjIGfvYQzhahn6
R/kDiYQr+9vlR1918mCyI0HomZOx7kk2rQD8/4UzKTpX/zlaYbENgXgEKC3hw4hy
GNUecpr7K8e019ttHWRX6h4zBDFOicf0JHDp8QfltvhT6E0ebclD0hMcRxjP7/lI
wHxJsdQQtF+bAmTMl3JuRX7+Lp3kmaMReK5gxfDwz8r2XWmaQQEowWOXlZDHuVt7
puFZSRbQNkfGz7Rh2aY9hNWYrWWJTYfaY1qUjD0NFyR9mZmLexnz9IS9k5QRqBj1
JGvVhWuA2asiZ5Jf1VMf3R1TVrq3W9ipuQS3BGG1m9cw3y4GHtkHW552ZDnurbCG
Ye0UKoZjusS+hZzBqbkaXnLmEg+FoOlcxS2inq6HgcuhEJbVz7hVsPu71glhAQqS
GXI12Ky901rG9nW8g7Nk28JuEYZzY4j682dYt8E/JOkLoNPmo0Rm+LD50heJstXS
lNqosqS1RhX7Ta/y9j0dhlYcMVZKEIQlS5daEk82TkayT+Nu/OU3iVX6UN0PwHWv
GiqvZTzcDUSx1Y0CLp4mJDAmtnjMLv7t12sgxKdSgv1AzHVlswKVpOyjzFc5li/j
HUiPFS2hX58KWHNadDpeA9utzJcYNWFjyQiTVOP2evi8hb8NTECYv83+KWbc0xoS
XJ0c4FxpNv6sToD269v4OsoCdh4nb4k8A7Vs9zkh/igTqI87SQX4JX9z0W+86X+8
vtawLVtKDWoFhA+Uqndl/rM4FOjWje6Ezt4PZBlfm6l4Vo5ivlUDNlvUKroGDo9Q
PE/pbJQn9dg3CxyuFSZjQt/e4HmL0fGTgBXE9dqPvPRYpjPmiCxdpGrtwnudnOeL
ln5ziFDOvShPwvLJ5HBYQ5iy4od3Vubxmvz2bsdhnM6vlb+A0FtheJ1h0oNJ7WdJ
PZafal8CpURFg9vJ9RTtb8BQuqFZohysvki9dfE+qg65dfKVSvoPITY0zfEj0JqF
TK4Hzvcl10o3XanIfVo+iFCiSd7M6A6RVOE1FazXS/4by8tuQHUy0Tqc4XFSw9eD
+pUSGufxtMEDb9Lx2zIO1Ri00RbGMtJ9N3se78S4isF+kfgbCfv/1IN1MoFlIal4
DuoIpY6vgbBBEF4Z4fNy9R026Tu1PBBdAtU26Ubpn2H3B0JIc7ea5+CBjpOoLfFA
rQmdgzqqVgtSWn+zjkxd/R1XNctGZyBYLu7ecx6HIEM7ackjpThXris1+sjol9Cc
GM4W56ThxU/Dlq/LU7rvF4bex8uW9nANXXkMrdm1SifvBUyd/o8WvIYBxebxdkDP
fF1azSqTbX/YKeS0Tx6gt2P1em/fYxwJtMcw8GI/DbFlj41Nl8+67zO+VKKw/AXo
hzkF2Q2HHa0ZM2GM2TjsSPk5QQDMVxc28Mk/CFJdbsC7zLLQ3rVgfJciEWDv0HBP
uVQY+M33VTKJ7UuR0AbIwxfhbbcB0fMZXDIoOjfbTsTZ/OFScx5BmWYeFClqmyvx
LAYL/746L7+B3QtzICtjZIURNb8WOAaLnHb60oFV60XOW/wOqVgrmHgVUkZcCwwv
AtUsa6uVDaN+XrtDsisKq1jyoMDVnprlsbxlmsbeIG/UxMPhJ0XTE3qF8/wV6xVf
E56s7daIjvh54fOk//wsCDymX27fg7xza+4aBt78azQx5jWpydlBxO5QwK4Fd+uG
0FuLhe9Cv/vjeQAqLQlbsv41qAhn12jGgMtFI6Hr6leLKBDjsFIb/VabK6707b6o
ZFID9JXYpLmNPdbPCsLUNvaWDLaQjA2FmJ+NtVa6ITOAsgovezpai3+ZR/LhrSUY
HozmEzwDNJzbsfb3lw6FfNR2LIDyTYolKj0r0iKklT7vEeZ5uO5U87m4Xfwlq/SE
khCcKI6rz9u1va8YLRPG0t3F3MGIsYCoscg+rT1oxgYM+4aeOGwDfSAbmvAeCpe6
ah3Uo/xgpwiyhPeS/IAf6yO+/IX5lW1C3FfX55phcbreynDTRvT9CTwrCDWbbfxL
5cKAegT8lLAeTm3EPiZvlogmpqryh8meO2I5qI8Kh7SlJ94PsRy+E2Flmd2pWymd
yQnUtcNOwcHYE1Wc1unHGzkVuxaFGO1eSMyD3IcVrVm7aMYJz9RM6dJ8Y2eCDuKR
3BkNYyv9oFNluQ7mrYWXFvMeSBPG8nxZQt6kv1haDB/fTgFzWcBvmA+ePl+8cFVX
I+tbaE1/80/OvN7H5OhI/NVKDyHYkx6GW73Yz9weQw1h2/As5CfLUA6eZvEG7323
o5ajI3iq/s+LgDEkRYtjhQ+zXcuTb+vuMrjACgqRc15HyErt0Tmv+mCUNst3GlO5
rMzz4Q6w6Hj3CvyXtwMuwC+NB51B2CqbsXY5A4l7Xup68q5aDv+3mUun6tFEOlIF
vzU52xsT45CU9E0PvgkgpNMuhA3A5g94lVY4fHQADFLV7Vmc2ALHKJF2OkCwxWiI
Qn347TZN8y3ECbX6qC9EI1BRHOEy1d1SCNETY5Kx+FdsOVfgx5tMe2J/0/BOUDIF
anjPd/KdZw+4DCxbUFsyxVtAqMJBDAsUJVEmZmBOZBbZfDnhTRVzs78/3k6XCxmY
1t7f+qPrBeF3ltBH4JukazgE74f519Js54eGBUlelxhlvGJ5w4gM39rVJH3bbZEZ
s0cx0tdSsgjMTSh9v3VLIATET8rQ9EOR0VvMmmIekjupM9If+t9wTPTkNRRk9JyK
HsjC0ChbR+lU6QpqTkwnjC+l4y1d+2QAoCI8EFmz3XgJEPjuh1b0t8qAsbxiNpxd
Msw0wSV4WY9nuxArNXuexQCE6Ma8emXYAoyNaiOvecEtOkd3jVTngFDCRiXdADN2
X5f9pqE95JBdkaHLmbap77dCc3lvUL0/w1a+ddxX1vWfudHGTcB4GHkxk/okJO0g
0cY8QBncAURPcc76jQzaDVXruBMo3KmCMiKtGuVXTi11ujV5hUOSWxonuPu6rBRK
X+bF2m86VvLaGv021LxVGwn8yvHexeO+HDAraWANkaAggU72SBuKBg7AmE3VoMuH
RJsupSg6X/T+QV9qyS7WqsjRUm5JaHGTTJ6FrWvurbP9z+H9RowDbv3aKTzsD5ZK
jjgIcZXCDyjgOVTb5bSqneTCO5dF4pIe4mZqRIjeDHUMobr7Kbqpt8em+FiapvOW
Nzxxqi4BeeFLWzGDAlQL3F7JHtP6MVXEWO32SV831BNtPormdoNjzN6nN84CEYZd
5dY8av5yCh5fj4gqBqfbblp7sQoc8C8aQg5IVm6O2OwtcaI4Y6Aux9Dqg+mTAjaq
yeykN2i37RfLUw8wp58tbpZpAvJorlsaxCzov93IfgZQ1bSRLLvFK47T5/jG2IBa
6aolhaZJZmXwa+E97bLifPu17T4Ul2mPc7qYey3Zt+F2dW0o8WeeKn3ouPDCMTJ8
fWGX43Nzrqg3Gld5pmwGrMlIksOZuSianuCoeFRj24iBII/Pw6KMJb9sxPOkHn44
BXnVe0vmIqVcRyI23L57U3kXG009i7KKwJwwmtzk9BFci/6JxpFuh68whYIcgkR3
41YhEOZ2gNoj+jBd0vMMYZdVQlPh5UO/48WBueeVYYFCkRoMuf9KaFQwuezYcjja
iYyCA/tTXyEwIvlRbBx5UepI8X1YUupF0VHlaXOFU7aQKh4GFzv/XcttGTMGPRwx
3s83x/Omisoqm98aINgDwYvo7JiAsUHJbdbIL9WvF6NtC3Cn+F9gBbKKGQUo6Kn/
O4zJ/yXAjz9Z24qsdrbrHfEydcCPuUM3DgCGZaITJp0Yx1N183BGkF9llNII/EMW
Ql+7Ldk0G0grbMMXm00k7dyeeBaSyd4adRKiFd2GSrIxegEDvX3QUPq+D4lG9sAG
lR2dKTaNAz0YbT5ehy+pwwrNHUI9hAr+lAVy6KYiJ9eojbyZijorUwQ5rWuZhxRN
l0OVVwsQBSXUGmuJGr+fLvZtd7X/vSr6VaGAx2H0CO5uFsSp6Fmg5p+MtN7SUe/U
QcdQaMeyUXqGB+8cPe2z45OlDWqF/WWFyjmJcucOFUMjM1TIx86gG9THRjJroT91
+9OgCHr+PDlMBgngJVzOYzTq62J8UZxZZSqgwY575vctaOp7SL2KUlJThsLJPJiR
eaiNpSEnHqfcIMTFxZwfD6X6sGGT+LRU1AUfjRQYoIJHZQ47QsbVLTI2QMRRJ3o/
b02cBUpohOmH4RdrdmMxng/xGwONtdh3h2P4DeGEf+dieI27QQ/GQhyPpxAX/RHW
fhgKmvSXox+xhbi+2WPWsY6+CVpDxQf7zzauY5u9F6kH8hzf4/tm8wkAXP3dq6bw
BTzhZ3UJIE31f8DP7vOL1Mxp4K+z4FyqX2ckDDDtyyfVttODK2xoXo5e/Ej2wrQH
2WV7re9BngM9r0UHii0hR2FsAl6BlvRgoDeY+vB8QuGzQPhbgFpMlh0/rSl04nqz
xijbyapOUrfRvsqvs5BDveV0/VGZt/jr1zxKeFI6Nb9sGVFOdtV/dbHC0tbJedF0
y8vde12rdMuThMCpCkCSnlQ+jo4viBZ4WVAFc0vh8s7ROVc8ioMsqk4mlubTjNVr
q19m/vA6npLHdfyJFFk/jEQ3X7gRmq5Ak+sOG26pnpDTvxXJvfJaWjXqDHAuzB/m
OcnsUhpo5f36z0mXvWrcfDBI7x2J50+OmjY8x4qSD6NsC+kO1U0Msm6MPoNvR21M
pvQUBG9wPeeHdLNU1sYJCtSIzwPEFQKCJhrut6asgEUdXTd4eLCj/DXtb1SUF6sw
CzsjuEkWtOYtB08tV7HWrBLJGUCgXxAiHDa8RYOW7qn8lYbcQDI4lWQ8ipuT2uu4
blPvpbysqjqePO1FQ+T/AmPDnm8OpV0ZzNMA6OsnZ1oDkKW9eXbhBNXkNQO7ID1O
AC/PMYQQo1BXAqhblm91r/pXm1Sq82ACMraBa0OzexwL+1hNv32oMYLaI2q/eZBX
EbTT9JVHRiyPomOwqdCnt7ZiIj+w8GERmRVwp7fpq/3r55QsUFYsEQk3sErf93r8
A4YcZbJN65a6ZqZfPYYOgvFhQUGUl8HO8wlz3FmdmDZD1ItHOQBONkG9E4oa8956
R3TjOagslnTbkT+hf0F1pOJwsVCF+fxE+WwMMeEQduzpNOoiql6s8bNc+sep+rGK
v+tq7Tg+ysz7O7C2qgM0al7nOFhyfWUwrrLElMf9lO7/8dVkTKzC1yeW01Rrr+jW
9E2uv8xFuG26KX7f1Jvko1QBWzBuyLSSRM6rM7t6qVVzLyLkobyskAXGg8di0w26
PlDuYFNCNfpibBLkBgrYodL91sYVay4a/oyyA5NMSfR7PyrjY0jolNw6hECqTP10
2YKJkCA/EVA8yThX/fD6NUi+UaBs3wVOfamAzWvFpaj6w+gV6ggabAcvLUs1jvlO
8LZUkgzLhjv3KEvbSF2fBK8ssh5NT4VzwHJwLB6XBhvx9SGGbUn+Dyc3n0nP/QWf
cVaCLFmGJRA7p4A8l8bQpvFKWuExBB1kyCGbw4XHMELzCCsk93zshQI/NsLOcj8r
HO4/5sSO26k6SPxmZllqtOZXWEBMQEjXIqBegsahlLbprSnMNZEWgKtq09fpF+3o
NOf3V5EX7iBG9MELzs8HVVFh4XykuuEGEj78MAQwvr36xU/SgG8N6uISqm8988Pu
Ix9v43FJ+E0WT9S8bgYIxAp56gN7cSO7qQxcgq9G9pjXrz7HvUiYBKqGGAXjIdfd
TCtTDpQF94cvJDPPJz5aEhJtohsyuq8+rtJx3I3Rqpcf/AXvIiHvcHlSuYY8+V5I
Lf0vWixx5YzX5E9trwLI3c02DAkQZY/02NQ1X/qZdkmBei1Kw9qNtyxx6Hk8sxCz
kxSrxcJM6pqhLzf92jxtaAGmK2c1IVhtRT09SEgIXTwmrDnpnPRQxcA5IoH8LdTn
cP3dorryWyBt+dSvLmB+mfdoAHrxq0USP42vyPyQsYDqUC75cdP4jeQMFr0hYWWY
ljyQIKk5tgzOWyvJT6TwpGy+mv1+mja/2f7sOUTaXGHVa3ysi0Jsvyn8SOGBlYOm
yLMqWm7jQaSpu2EYdhWojM9DIuMW8b07doltxpe0hp4NXxTWq7VsMptvUxPwAUVd
XIfJ8gCiUDk9PgC4YHjiX0BpivJMBx6xt7IB7R7VywXXw7T7wgPeOzD9iCmflK93
oaj+lfvVIe5yXkWI0ZCtGm0LHe+CHnGzFaOcEah25YPO/b00be8nB5D3z4DyL+ll
13IMljRUzxCcCHDx6X61yZKIlYqcL7MvtALC+jUZY/LXFVh9CqKirR+UTLaZjVBu
qIk1wyow398nMVA0CH/TgSogExeBwlQyOIVTqczTyMp8TEjz01RSd9iAUQBWEFGN
YlaWxTswwK5l0re2XXmDOuiNGSeSnLTWrrhW6CrcmUcCkdvBAUqb5xVqj/lI3WvW
JmQu76XRGshcRD717tswRTP3rHEERMkgX2/D+Mrbn+oI7ePtfYr3ICgbwQOMurA2
7X/988ID4pZgAmgz0MrcyrRLs4vTcCL7lAQ3pX44zACF4yg0ZUtkZqEb4tIDBasy
G0Kw0UJ2k8q2u6olf2eeTNLdyuk6RDf+LcPnywXx5CvA1tQfiiV5dy22ydQWIAJx
dMvkV264poE8Lx4WVJPSlnkYcIGM7Dke1NAuAhXWJb6dOe3HSvtp3DpQEO9hwFe1
q8laot2Ea6BgyoaftC9SoSK5RFXT7y+kNanP3JttL9rj+trcVuHpuI5e1gL0SAau
i82LD0ZfcgI8qefmPCPueFlvcEhW9EgfUPqZ+p8Vbpmu1APBzyNxPsV4CFH0ekcL
w7lPU6EoExnZ8FDuu+cLzNTMWZ3Kk87zL0Z5ZSG+29w0wspSk2ALEm+uX3UdkCdi
6EuDOPVDQsUKrIsqIIrZy5IzzeaIQATpecgUlfXNLkc+tr5WrxDhwoY50mFDzOWE
zxhoJHNKS8+fHBESaoTm8y506t//FGri7BbNAwZAIGMX78dBlX4Huvu8pkcVetYO
O3r+mAxzP54BaIRBy/3ObwJts2ugmsqbC/7MvfQfp3As8s3dspu+263BL3cr4NSZ
b5SnY7xjpG8hPg153BlSj1Lv9v7d/SI1IlFKd1wEQoWrAQbz+Ue7rH9x5eCrBe8E
NqGSMBCtRNfelMl2/83pNII8IVYevo9sIiLghzJs+2J3A2/GGtd4LtqKaW+tJHbn
Q317qNuEc6MI1ADVeoTor9PkAdftHIJbWen4VdS/hDZhtwqOUjp9zb4d1LMUfsaA
SpMMTrj1wZdSoYlJ339jmIP4EtNUvMirbBIIRmeJwLkzhDUL15lwZyJgHaL8YHa4
Xkt6XaKfRntVAE/fpeA3xnItatjovP0KDYvmdfrk4k7DPO3jMZdFukr5VX7WO206
6P2D+jSsLwbfWllqLDKJpqeoOX7UCAmfrm5UK7HvK60V2P4qZlyQsv4vRCJGx2TA
TT7jgAOYFIqBEWqjB+goL2KOnQF1jrnRklBH7ckdruK7LhxTgbuQZiFL3MXLlZOg
d72YEmrjRbQXoouTIDYPcuJA2JZFZCTSbzD6jIvPmJUThZGq4N9O46B/xkII+dFe
hmKTwfXjswa2cyRyghkXzlWFsmhwYrJnA+2HxQwYQbe8kNAMwBc4mEHiRlBdvg/d
LowG7TsNWZJ3i479gMnbfIXDWD274jv5WSHjLw5RO3t1S+r2AQHnabXfbuMRwgGc
EMDvWd+XQfMCGbbKgXsdNytabrMcEXZHHKsupdlP/rvPPYMhdpaisaNXiArBPCpT
gDnkrQI1Slt2bBmicwpDagTf/6qXaC3vIht5ieh5TZdTL8YGDPkQU4mKFd9VNZrc
sZyS9VH9iQfECfE5v6tAFfmP54Gb9BDRjkjO3OaeEAb93C99MCnfWP2M5rYuAIq0
3BHKIELTew2xDOkjoAg3u0Ai66JCqXHuAEE22rO+znU4uQVnZCR4lZZiRSSbCDGf
23GOS9Xeod8mFhZ4kYtD7iWfRcW3ioeEwFSqQrlkGoD6RXuyTJ6nEnqjYolTNs4q
teLO3n98L/radv5Lo18BVVTbMeUPfgMTgssF6cRTQ194ixQAPtbTvDyBtpG9vQYO
C0iSqqLLY8BfcuNiICK/S/rXk/p4r9FRetNEdJZsQoel4fxh7GJ+thMpdHF8LQbO
0CpwQLdWgpL1y8Flu6Ivur1SmQUTOiyWNz5jgxLUn6XF9hMjCjCJDH9GaVglgJib
84tihYxx1yGefrlIz0q/BOZ8Tl2n1lHyGscKAEXsU4JJUrE5DtvQKIkygAdOzr0/
5rKepkmPZZONj3y/pI7SHjerfxwYNQ7x+BgblJk3j3T7XIk2vZgr+wBOTaFFZ0gX
rCHbWKhkAunNOXoChWkuHTRQDGlG+UyD9eb7wGJESyVcKvWoOiOHq3LgOLLo7ueV
xBJfncqsItocO8vSM1ajse2ZDeNt/TKL1YZNB9qWrhJ20d4X1kWSBl+7lln+aGso
uArbmD0xuq4uQsRLzHzavNxZCVu0dWR5EeG43kE7w4cVEhIp9QBCgfJyawtUatZc
L/Mp/oXH3nNlyHXreIvSyrR0knq/J3dNQ34ByO5FigIZEmn2zc5Agu8bjVgn7HVL
morYOcQRxkxyDerywsjKI7YQAbivKfPgJIEwoXWTpuMEtMtz6JnrHepOaNHFmx7j
nAC6SC+SuGgBPHkzqcaXuOV7FHK2ZKEUb9OO6JQxyTCBIIKPxziIVYSRC3Rt7jqN
QDk7PTcM8Yn1M1TfDr/0c9FIkuvQQYXa/zEGPOi9NAcUjkhXBEDyT8l4ofhrJiff
HhBz4RURu1nJ1CjxkiQvqraFcslIAUHrm9bF1/RtaOJelHxVxt/3pNfqA9YqSoZz
qGBkIEQKa1vhsA4ZVf91waf22ZhF0UBCYLoAfs1LIUru59yQGOoEo/4UTQJixdWi
PHUWziA2zOX/KliVjMcxqkp10mwm0cdt79e7kO1RstpbytUHW7xuATbdPQfuknPx
lo9GdAj8zN5pnKo3FmzwqOvQMsQXNKx00ExxUsHtPwa4GYrOtW1yyd1i2z5fc8Ac
bGG8AFkES94cbuf3OCd2hTqH/nqbmCbBc8EK2D3Yc39eVi/bZ3XWsF5hZblVcE3a
NAz0PxawDv1Ly5loDONPPteB6bjB4rrqkfgCgz6W+NPF+Pfftj+Xdicf9/R+UtoU
0x2htmfH4waN8yUwLW7ABq/NAONhtX6LOqTw4gAogKpPA64Ic3EwL5ph5CiMETJk
cw+62HAtrzvfAjSxtQb/kF9tcne9SaMiw0gISnsrwxxucQ9X8spJxSEvvvwFo8nr
zikIYZUzQ6Fbya3P4Zfjjy6Xo2cX26G50hIF/ZnN9jW3auPaX4HbltA/tDpqrDbd
v28CEUNyt7pAOU0Pt8LgPw+o9mo9IDlo7dTnU/BGZ9Z7ACjv/Ze3x431TgVGVxEo
Ej7u+bRTFqXnC1MdC69qiR8tYRJvqBv+JWSjO3ZkXcB4ZQ3z+Kh5RnzzmKyH1AHy
x0xMgC4FUVEQZfBDL8ko6RZaS/u3ePI9qHXaUIw7fCU+tIMXLY2f/bk0+tQqE67W
vL2FjMKGUhmZzS7+gdbAPs9R1qIxzi0deATUWGzIXl6b61CFdUmYNYEvILJDdPp7
Cuv5dH2lLCtcEIJuAjs2O0WPv2Rf+lDapRS/jjdHVqGwojSvlUfQKu1kR8sD9YCA
Lphf4X+t7iJ6sFMonFRWTlCuFycq5baKZd8CGnB7Wy9za/zAD4IJj5fQzjH/F6Zt
V5pOxw4H4v4/Y9N34cTu6DyZn07EYkBB3TmDs+Cv9Nztv4o8HssihilUPYviPf9/
86oJGaZVoG6/CtgNVPKZ0MlvxGzXdweKqNuH50XdrnMJCow/cgP97VpnDQs4/TBp
TUDzArDjF58gnZ/YS0l+lU+/efeNPVJPtHIaM0AOXxy7t7MhoBcv4rc+EzRzgYRu
dwrxeL1Dgtf37anCsSdaVOQM9b/T/HYc1xUG3M7LJ1OS8oB/XKCvMEwceuh/efZk
0fXKHadMcEQoKYVEufI0Ihmblr4zSgKzdv7QVziqLmGtU0tF+Ar2Ahs3heiYHQrT
MgOtZJqcH6x45e17g5mfJokbqtKjyyDRPNmN29sgEogU1i3j+Tc77T+xtEjcanma
jG74REXlUJcD59OtyPvk3IuW6FZP4ktZ9Ys7f0f5xYZdT+FKsHFMGuk9BMJje15h
nNwKDcVRXFQ1yeGnPjhz9ar9O0izZoyM5+iWYvII7NTmlYM77rKDl9RfUBqhejjT
+E4MNzbXiKzMsbAMm0drCfOIFTP6RJ+ImUj/hNpGSKXyzNfyIsoiZZd8gg3QZJZX
pQHv9vhrkVUE7IP2qQiZP2HkpfDtLfJXdg3CWPDaaF55B9NJgLttMqNNHUH3mCA1
hJMK374HLGATapUCnZHa8l6jVeUOBcC9aO4MXnGeB48/9dCXaLkx+4T0plXGtm1t
BLZ+uM2G2QPtTAiLbuKe5fQEwSw5WX4rvkb6XEXCLZHNvUNHQan3LxZf7zDwvPbS
fgUqS4vWdAKC/0cg8m71ZKqBi8SbF0PwxXXUU8qTmAi9ah0FFI5sIdNK5z4vvjnA
T7eEhQohGv6d2Ta0F2UVorT7JNLV/MCMn9ODRhdsjSjkqPiyHnXLvd0kphuq3gCR
UFZi7QPS+SfUXJpXNNW4z+PMEv/GBMTXaY+ys6GZZZwYxpm6bRN8N1MjVi0FOjsW
00r1e+Wm6q0MVfDlLd9zy0crUdtKeAu95YxFUhnMuSHGB4Cn2cdYbX2de4Bt4H37
r8+DUSRwLSo9ez0kAaM/T/ZQLifg34LTrvWdkWCZvSqlbDLASx5CRnNE9v3e73jM
bhqghzLo1PmGBEFRpjaic9kTetoGs7PYOkLRqXmvgtFZW49K0zzd6xLhfDRcnBIu
GWE1welw4Targu9uXe3ZxOfvooxMwXpQLPQDfFNrdD4oEMTKN/B0+uzW4Eq8lEZo
6etHNK9swtxuq5PU+qUifg0NxElxfLJF5oPX7WK3vl7LFJmgeKkrt56rK9K2a82e
ExRkO7yEKMy0qwAAiqvBiy8k1rhAYNxS0a2ZmcfmjdZD9YF3IAkPHyOU4XS8dHsw
d2Pu0q7fXvVJLxmG2z8bA8iGmemSQgp+bYkmRxGpYIXBN8bl8c6M+Wq43gmkpArf
TiyI6J2/0DYfH1HUvU6KY4izDJs0sNev/5dmH4wJNm2vXV8YXWj3fpx6uwVyQqix
fIxLfQ2Q8qB6HyI3z4Kh5HVmhZhEi8VV3LnyjyI50feHU+7/MLFfIrQ0Z4Z+ogY6
n1gf+HgX7AKKQ0qgPKrWxSr+NNCycCm03hTWmh/bf36D6c2KubhHMV+/cCBRhJo2
bKY3Bd+LRXMS12PaUXeUQ7n5UPDYmoYXMqgEo1adMjnch0Jo9uDejygpPql7oEM8
l62rn7sTbIzPVwmcSJpXHM6QztN7FYUPHvQBKfHSw1NvigZP4nDZKMji7t/rQsMc
nK8im/xVkEUlljc708bzgXM/lPlV6SY4ixURyyIsc/RJ8UL/u6jGXv456vPeb5tx
1oX3oGKohAB0sEkD/1mA/cQZogETf5ehHKbTatkdmIVmL4VVs9l4dY95DJuSzr63
FrVaLjouCaPZUJf0aw8WUiUw9wCYYYk1cnUumfIht7Zz6OiVUStBvonB4KXYahYe
k/HzecdxX0eCVJRLGyZUOPTtPQSsplgskRKLe272MDkXkGuaCtTrE/q6Z1eD9go6
K9zYg+OaDjDMQvPyq2Gcu/oXFMvxO1pz3L1hsNBloje8O2vJwHVv3UcGhyO4BZKS
P6SOZGDyI52F4I7OquwGYBkNCvgAOF/TdbWhfJJwZzfeVauOnws/U2brp3nKcKBk
2HJLaakgNvC3apU2/ssipMaqE++jV7SfuDKz14IEDxUh6N8NSpLs8/yVXjf/jiC5
PBSGAL4Ik7yqXEBQoyHaP79FNlmeKhCbjcG0o4SpwRHi61LVqt8iW0YHoRFier3D
HgVEvDkgFtlE1RJIAR1v0xE1ij9fyBeVxMp2oK02svhLeHKLYiFPbPaIj4san44e
vMRgJxPB5apkWCfOzMqYpFRBvdQJ5yhSW25s7+82hPqkkO3UTQ9EOJT5Xfi5H9gu
g0hqt+qSBfnlYqAP4K+FdWBM5oRt6L3qi/KbvNXoMFMY6PjXiSxEENuKl7b8GTyY
yT49WjxDcw5bnPAcOvCYMN4vzOK+h/UHaCypNMN89sJO6i4HYkCzA2mrlqUK1sOV
CDbcovJ1hAAq37k8H7FETCrRRKRew2FTqBIXD8q0B+RRkoUsWBgyWcOwUvtDkdkU
ETnzvpUyI2gApySizUt4TYnjGlW5Kikkrqs16pD6jItq9IimJhvzqo3R/PZpGZ4y
XonG43Q1pwNkqK7rHl0oKICHRjuuNH/JYCIN9HvOA7DXLH8Gwk+T8ZcHT8Boz8ip
/P0e6KIwotFV6d7evgxkfCbfLQaQUpRan6QKyKLPwEURNmX4Wbu0onnnwVPlqmm2
MDD9AV2M8ujmGospaj9zc8GIpD2uRF2L3/hwfKE6+DVjy3rwJwhlVDBiQ790jW1r
RVlMZ2ZYy9uKZ3ZBqy2NFnG/RwvOIRIJdfBrN1Ax4FD+NF1F/VzNQcTqiaqrtVnR
pC+J+nLQjKgY7pxuU1Kc+yU7n6PEJsh6qWPTaGibSm2m8j2rVBsXKy5s8Aflkmyc
mcDcEkEirvzmUqb0HiNBapKTyNqVyDEkBR2AgVKVkgfgF0rp8TXsubgP+Vfc5oKQ
vzv6KdUdsGj5I4oj+kPVBSDBLT0lr4E9uRAMTnsS5XSaUFRx3ovcmpai+ABg07Gu
8s/csu8Q3Lk0yeOzD2/OjXPHM/paF3jadf8y+Jbsrn7JJmRb10QWlvmSIPD+tC/f
fRaAcEP7RpNGWbyF8speh1bC1LxS/b3DGjs/djVzswWM/zDzJpB1ic/z21N/R38Q
dK8b5YkmSwCyuROz/o8IpVNrQ3KppUwFbZ9buw1JI20d+d4jis2m3BNgN/SDZ7+2
HzBG/DudOuUSZIrFH0qwZHROLqV7XzhjnG158wM48czGoIMX1URFreQUSotMhmux
oFgs3ulMEBvMGnSEFteGegVcWXQLZX2X8OwfWE+NhriZWKvyy9gMeJhDU7wom9Eh
Tna13G6Z8XyYD3xMy+5ODDw5yW9Sj8vW3hY5ON4BdzLZh/4K2MVqXqD2FQ73mxeu
BPWHn91r6c5t6uXKEIn+9aAFoXZLQOYk2YjdXBXCy1SekA3JnUnXxBhAtmIDXgrF
UGmubv3sj3z01ZfEy1t5/FRWFGASucwwCjVdU5yLwH8lE3muVy0moBM5AfCyVNEX
fvqsRczEtQ583b3CeKyO/Y+GxwMMHA2LSHzpfNrAnom0MRqYGJjHMk8/+hmGDEBP
Osp43udrDBxm5QPvpKH5jWkvEz0ZauRAPLKJuZqUZ/tUrtJ07PlbVMXQ9LXNI4u+
8xofv/n46R10e8yty0ik0/DqbqYYCaTq9qjsV8QQpNJLb6RvJG14kgP0m7CsnDVa
x5JMWD4oX46p9aLD0AuTFqa2uGzdrV6ILfCwHmRSUiNnmWjIU1dyUCqUF7r6J6DZ
maVR52ELHRLaCO5A5qL6ntlp5MPjwsnc1j0NGEwMwSLglmaaDXqOXLLgtRTtmhf5
UyDonc6ALblsZJXFoExqLtCPreC7BJ4jcqF+1s0mIdseJMlmf5gQm9RbPfhZszz0
LlYQVhWWrTcHf8xYKOVIR/XwfKBVtaUderVZDbDHBP1IQMrtHOOt0NZVjPFaZcrH
1//C5oXKPk7R3d5k+TljxCUONf24G1XQVkbYCz6JxvDIJRFDxUnQ255//YRjwcwv
N9Jv8jPFG6ZP5uy9uVrAKD0Ig5bjvNDmfwRxNpRtWQzBvuDY87FIL1ic1OK8kAZo
xtErVEaeHyud2YoL3CvIr4PqUMJTD6NiYKv5mYpyi+iyrkObyfAnGFnntMZBI0Da
iVv6+DCN4pmsWzEMcf9V2FnQPo3orWgDNd12L8P0FFxyy+mG/w0jParyD9SNWDPb
DleQBtna6BZVwqGwUTG2+xWossLkRLT0Bn5xgvrBGhJIDXOM2kKy2FGKBnPB8tt2
i/DCTKtFzWvBoI0R467+zqdr1Mu0eBj9V16QfFLd3pf4R+wowSC+Q4yjsP2QqLj1
oWSg7pv4jXa24N0nMAg5wkkE9uI7vIqkiZb8XxP/fZa2u6YQNYOI6GJmE+TfdFzT
G1f63i3KyIHWFF9itMHztg06odJFsp5oCNzpCYLQlf/Jc9/whpHnQSPupwk8BvuN
hW5eY5ucjg+PnUVi3xKQpTvUkFY3KrlF3rzjYonZqmInd5qyElJ4zmb/1G5NQ2iM
bc8Jwg3DUwyZf/a+ik4AkEZFC7Sy+eP4dno1jwcHAuvSy/4M9XMWqKft55Pudhnc
eITrPC48aDV8PH85jx3+17YZCg7syiwNf2nj6XH+BEBYpy81/xrzqShiLJHmlEl0
/ro1XwRiGJEIhUoE0S6jFU0P38mEqWamTVMnZ84wHt0siwDIpv5lXX12i8+GL1Bp
IiGu9JI2j/t9Sm0haIvE2awG0qWGITPawdK/eups0AXWrD8FUyrgtS731pzluuwo
XRjxMRk/YQJB1niTtj3Q8t+SWTWCeAPtoGPxzQkMcIyM58B0EnrBqilJFNhvWwPY
a+siJpTFCDR/R3m8DRQTrjwlrtyOUjmvmyF7XUSibRODWCy5UaaVQr8+yaAXYwtY
XiSXVu5qxDc8QF7scEgj4CTg/BPxqwr3lSLrfH84K9moIf5kW3unkIC3sJkmSs5y
GJVqPmYeBve/ZXosRWgaX7Ch+ECRxysTaJ/zSLTi4wTBuQjl2nNkKgH1uNBt+qiJ
3xSbmVGIrBT3ckfEkr+IbdE60I1TV7RwzBIFb19EPZPhD6+UO+FQO58eVoluQzXa
WO6XdP2nqlUbje3PqD9AYZ+eUNuaalnDsscMqX5KTa+GnzoZoMZHrXzFEBFo61vd
0gDIKxyPhNxD0+6zlbCEtlne4sphTMwMqMS/mxzE5l+yX/Mb1biU7MAaEwDafn57
TonTVbRB1mBaAJU2Q4izgWaq5qHzuIwP/APfnnW8m2s5GDidcht+vmY+e/MD46QZ
+LmCIvhw2H32QGR3itDGgXallwixzCq0l1iZlTw9z9sYYRtyBuTgMa76jaj0vQat
PvF2rQbSuaHv8MbBPj/OlC14xUunIM/ZItslE4lLOvLUHgTgR9UzT4+2PE6gzJ4c
idP2bPC2uH0SUbupWsjA5+Czk2L8gqOAtY03hfvbZOQN5sVzVd8PyL/jhM/VxfQl
Vs21rRH+RBFoEHaxqcbUN8mS1pRzE/mW3iW1tJ0K9O8xr+8vhICv+Ek7xwr7o1p9
KqM0Tdjv5eh8KK0czxC+8EmCkdxWUdx1eI+UT6lieKPaS5CqXAC62nR57Q5Vu1Zz
F4av+IlRjDyikRluFgMRGAfojd1qnKGrkyBuABkiX5EUPjApCeVxGQYPTZJ6IEwP
scr8dE3QS0ylUgrTB58+ZQSh5rk2ODvvYDgh3w0TdvCCOt+LvrVm3RQUHhNPJyUT
0b2Oi0RtqESLDHTktloKBrZbmbauk8B7+EVt97Ju5iD6Na3gcgmxYe5aq11yPsC9
FkzQNhBiwwD34oGZYLV3eHZ02IQPxhyLlWbcn8RiE2Q2jyyREr2CRcHshgWensZk
suTSG1b8voE0jDehcuBmr0t8pn2+ItWi5CkOmqLOgUQ0h9MdZr5EhAxv9A33sqYy
V4Gh7Hq0/4zGCbbiVl6Yp+ufblGJbPWObQNr0s/BZeUKQf1ogwLWEvRX1VwFzlc7
+72ZUmAL0stLtZo3SRJL0KgispPFrDFNPoPOu7rRcDFBPOmwhx1fZbhheg2JmVCe
E+drQVVlOLX4oHXedb4JWVtUFUsa0NnfgkmiJTsm0hBmBVLRl2tzjYPW64QOZbxA
t43tS1ZdNX8UvBzwR/5UArPP47n4s7OfDoZGqJkTrE36TNYfVlSMsMYkvjM9f7+V
cZgLLQkeickA5kADBrHKgMaPrwQ2taYmiCWjYF5WC6ubz46rxPf+1/5hjuH0e4LQ
WiRDdNxlboXcuSTv9qCq1n61z0cZF17HOuGdQAjJW5Cads0dlKaOaeHs/QcqCPtX
qajRNfsfO4d3qS3CI8L4FXq6ORetqw1tD55+5mZrDwWIMKWuVov6nbL0hKOMR1kZ
9v7sVEhaShnW6CB9m9FXpswYU3ZYXK3Xlh7OZtuT0SHSNTn8WULlH53ZKkjyawi/
EEFwkmCHd4+XMYbJc1wJlGtJvDB1Kpi0JjWOk3vCJwO8C9wGF8Hu4TPoaU6oj0Cr
70D1KUslyJFsbZ6HjYYzKjkFCZL7kzMXdSRCk0lvZ5fzhOu/XFDJi68nwlqoGHqs
EoJ656BPDa88mvD8wNQSHYIFfRQIz4L3wfo1DgEqkFFut1ZXZbFCfGPvyMJnKSJi
Rkmy1fCkwtnWTxi0MaYzCqjvy8ljZ01C/6QILj8hZp6F444XfKDpeNS+25SVyqNA
Gb53ZKIwQh78rz6FMFtdMBVarQm1XIJRoVmm5WxBs6k4U8mev+O1jhYaDXhuCBX9
uSQT+XxfwbyD4XgADem1t7aRGjpWTu0fF8nCkil61mfO0+G70rmjYL4HeIKqsihA
9PqhjozD4gC0iiPhRELW7E1lUopMqyT8ArjgrR+qxn+uwPodcE0zMlvC3pgK1gvQ
Ex/YnixLrGKZX8uEBg1IBothqHyErj5O/HBt6oTu48udBiZ4QeXtkjyvANVVZ34R
s4GE/9dRr+ugrFFNJSG51ubSdrKaIxa8wd3BEgbJNzI8lrmCYcWFg29oVJ0Kr2VS
AVi+FSQSCAbxwZDGowzX0+/BEgpwobVywH+Pjw1sVis3AhwtkA55relfnWcS5I+l
N26DLKsj6v+0VFRiSfG1uV5FKKNcS9COkgypyNiyqgO7eNZlUx3tZhgagxyvOZmo
GYgnNjXu6auJ01BVQlcbQ7aPO8pAchM3bb6ebzEVSo3fLi5pLJOOYzpTUgvxAvL+
nolMuEpW14SJOTomjV4H4fxYcX09D+MRRKDomcekWZKE7ae+dKVFtZI++pATTraF
37nsi+pGZrXTwmp0aSx08FV/cH0eWue5J9szlgQBKQrnzZloUPskP40Gtyz5fHYi
nm+Fms5wj0uYN8hNQkqSMczcYU5FradtSVJUQ8cCfZOUONb2W8kAnADF0xLQlDzM
qJebxIPZ5QYN6HvEsx07kgugikp+zSegWdd6Eu5KAd6vWGKdxuTuB97w8K41yoq6
auexz54gpx/w4Nlg8xwShQrXIIaxEVG32KAsqz/HfRowWmV1nv/TPJ9w77BpcrAY
AxeO9iGdnS+e1QCEd2YuvZeZa9yh8OBWtDuPZ+y3IQOiT9rQ9cSnmf9M80PsX+Hr
xQ/MIlE99CHXkyEoeoNhAqyo6SsSja2UStHLqJPKLsZHG+/bFC/XDq1IWmoj0WTP
ZX4096IpNRjjBFCPfDufi9tx4zApHVDPnZLFKXPDEs1fx4Dy1hDuz67mD8TlBnD1
cNkSTQ2ar7TWFDoXIe/oXqN/v46vbfE10nQVAh119wc8PF1zGysoNmhMapUBMnXy
fkf8NX6GRhFUsb4iQytxI6ve1KHYbg5kf19COddEn4gmjN9/2Jl/nhqcNMQqrjRH
NzVdzGdTTh6i5sgNb5dxzURdN80iTB4dpQxqfRl3r3p0vt1qSJ1ZKQe8S81aP3N6
P2hYpJYpdwFt/Xt0tYbRKlwYX00PrYQb1JuBXWEa7A4xUVBdi3jgy0V4uTb9b31p
+P0DRPqGJ8GBZDH/r98mfkydXqvJHLiSF+eh6TycxEaIehOBlirgSUJPwzpl5tX9
8ZcKSqCLMUjBMHL3myb1nWLZeL1WUWrbkkLKw8eBaqfLT7Ip9HOJljnhVL7FOpYf
oR9+Ohh4qB+INBcOr6dLbeAVqsvtxvh8SblCcL0g8w/69gbRByORHM35ELdovwoa
2ojZBItC/aazy8d8jklhe4fmBPxzkHjXtxjtOqT09ojvTCvZnElEIfnX+4W9MQuF
srf+b+Ev1OPGKlbXtFlwg0RM2tJ4xcgwMwmIuQdOOmO9tyjaT/F+KSEbexXTZTia
PXcYpBP385RH6LkfQKP+IqWjtRvNVb1qGm6Q5eaICWm5jVRtTccZ1MhloPEAFHbM
Ud/yxt5WK+RsqImStSPr0fCOdO8cr5Y58sRXv/P93M8gKfQEFFvfxM/vZ997/k+E
pWUoCGhlrLWs5mjUv+M18eYObNMZ4wa+1MX23eGXXkeoAlrSAVRqLZuV4pjLhpSR
FAE4fj7LgsnCOLdyj1ltFP54gU51la8BSHTrbcHdaHVFWGU7auftzutHs12Oyeov
HozLdya70+ZD9l2vKo7UmA9nyiaz6u7AwpqKM08vOjFIEWITLRO6QeIktzCjLs5w
BtkpxqcBFRjCop210MDZGSASiUBScP0YVQ5KjvXAPLGgWhSeN9KSHmEJe6Mbo3UU
xmGdYXKSPi6z9fW1Stid+0CG9s8thzHL85wVdyxsBkxMWNr/JbQKW7s69QYTVYaE
b/9k60aMZq1484RAQW2TKgjffshZqpj4UCGOdBbVNxHa3pIzseMt5jJQ5iFOZWbj
GlEqlKbCqoa0c0mJ/hvqBVDcJCSLUzFCkgfafsatRdRWJTlQZqQl13A/G50dM/9s
xse4/gXMvGnpJPHeDpJgfWsIGAwy41XNQunTqWvHBPmH5S5OAr2zlYuiWWRgby2V
z3NV2DvXCw3lm0VyBEZMrsPUfWm9rd+UvAmCycwGkeEqmjPG5cLm1Fvd1Bhr2vES
7de/4lHBpblad46i10TFysXgJ1UwhigM/CEDv91BjmOd422emyFMjNklwDAlOKtG
4MkXf47jEH4DNrH2FYBa9rcKCV5j6/BIrNWWZGuxM3inRVkLNspx4Rr8CaTAQ4wG
D2qk3thCiWsDjFzdtwW0vZ+Lxqu8VZlozWJ1ah1tnToKP0dk9GSNLCIft6xp+E5C
qZvi1U/68wYCbvJ1456waKcXteTv30TIE4SOaqFgFIwfIZkHgD24i9Otp8IBDKVu
9VKMGRFNZrsRCisP8Pxl/tdffWa2+JsiACNbgx95L6qpxosi3uTgIEea4ffjPwsG
2RNHGluw2HTicoG0Tx9xB0TS98Bux0QDimINfE8DdYSuZ9P/TxisAGhBArX+bSj9
sRuHhs8ENgTbq+tWH8CJlHxyoaPOxF3pWZ8ptWB8+pc/nTLCXEZkO/hqtSSleUlv
uBBT66FPKz325ga4/M/qcoF2huhDtSn94TEVjhnvkRxwUmKoDpKIipaCF4JYoJLF
ZQRGI8AASLnDFyq+OARDG6hhcXCalh7DlUpxZiD9ZhJAavsRhmehbkpEUp5CQT8T
vQYfiDJ1qHWkboGIMLwjBhFE9X5SblZ2sU0CcnHkEDe/tptHDVhhVn7KmgH4l5cu
5yOzPjNypAIS3EoZ81Fks9Xsw+V3mRZHIOgCDsVi9D443ddBTypGP6h4A0v3dxlr
MFPR6NW5Fzu8BWaUgbpAqIcrQZcH15GvED13Lym2+AeXN04jucqkf1cKKTamNc3i
zgGSz4vW+/ZIKSVI2UqAPYmnVR7Kvlzg2fRPwqZORid5nVS4XxAS6pTYbjbDrC91
JK9TwicQgiJyoJQuxA8xNYoZGga2Wuk/qYQCqewFkFPpaLciFPHHfwKhqclFULTl
4hGgb1G7J96eGKVztcvok08yPVLW3NXprDE7bgEvLkcykVdjmin1OIs67vc3AShh
rVE9Cpsx30jnEnZ9PqiHOBn9weIffBS/sLTSLJGXUP0UQhaHzzJqDw4EHr54Jbv4
bJyuc4k/QHHpTLP36EhOLOM6xIalyoqTpLUuvZWch/o0cw5RQ/H0gOxTFE9Poa0L
QxKHNthgRXKRgHHd3JbpSu2q+i+2rTBGlPN9+JhP9nezw9pEzZeyTjPvQDxlVH05
weXc3bNAIy1CnkHpc4ySG8TU3wqtOy8fLIPpx1ZeYrnKiXMTQZOA7/rK50UpRh/q
vrA94vuETMOaFw3j0TZAhh58/tFTwiTmKCMWxEc2gqnzb7HiOgyCYesYOQ1BiBZv
/4fZsxmZlmEZZb45MJb55FQkumLQgAiRppkpnG3PEhj4sc8QHGZYqjvBrXN+86lm
ioUiHMMTHKXmLvJVvMGyEfE5MQHq2iwN0NaKmWNxvFHL+5HzNPdWfTjaHvafBxhm
TwusJYq+G0sBtZfSk8E36mZVv5OuPhdQmJqzhFPrIV84Mm4wxfrxMPtp7VTDWwQ4
OnodPDRlysyny459NKoc1pPxyE1kVMpvSs8tfHC7Q5V3/YLn4PE+qQuiQv84lkqh
rgNgphiRSEQUvcbp64jxmgTCq6ZWXJ/AhkrLvAWZHCf8r3JRaFfdnKo2O7TseN+V
2t6WGTXKOxK2m7/q1T86h85TytZYcvnhv2T0nKfQTW+p0mPdreelRbQmiaHx131g
CY4b3n4s2MIXbYC4G7sRgrpIz5sQVvOHhyzEHRHtd69SgtxHXbCG6BgROzC5pQxI
W3me5nFklvECrVJyLQip/LfARXWSIie3WUzc+DkAR5KWjnmykZ1tQT90i4kUC/X9
kQk0dRNU6XKnSJc+ag/B3RzibSzbjCKKABLHxtz9jUmJjEYISOWMj6Ewc1HNu1Hr
pbmvo5hEbm6aymDrbe+TBFEqziCUq+hBK/fQVDgyEdW5Shyu1EEXvrkOkEZb5/0/
UzHwWPD2qkQKQloLA5JePd2V9hcWoFfiFEUs25tLUogMIXNoarx9OWehRFCb8k7K
mF7GvuYjx1rD7wObSzbtb7C9U3LmkIDhPduGSZaokAqR5T/jPTbJ58ljRQxB05B4
rdmEKUGHu1gRjRf0bo3cFJPwxRitAMY/MIQ04C8oTZAR8X6k8NyGAysqfWwhLAzO
Xy3xccChcmVzg6mKgy2OcSi8rglANGwnxUuCwRF8I4j+tXlppF65jO6zogohlBN8
WRLz//QZJKLhe71XYPAVqcJYKDyX+uoclILddZaYSzavUGrt9/4nZkSnCNbhi/qn
hceaWXOzDHmm/LazPzjP104snabL6Hc53DMimM9yiCn/dHzeJundGBNrQBR7grWd
2KxYF1pIjk58p0Mou48hX0/DiVYOpQbsuPYq3jUOf6yhxvSmxSYgZj7o9oh3j7+K
o4vtgswHjg0v+2AbgBZdYPsJiK+iuFLSeEg4pMa1eGwYrlBtjdt+PKwvNg4X8YMu
RYyZo6s5E2BTMhwe3H1WvU9dKpE2e0L7MolpPD57quvKlCK9Jf6kFAIJWFTg7Ewe
U2On0dgkGNOll+3N/h/4zs9nje6M5M4K4idBu9xmgK54dMx89kYx8nKhGEixM+My
7iFLteYyp6f2aI9DdTocG67M1SI0eoJYN3BWpVDY38t+Ciw4sw6xDX55kdb6TZvJ
GhRYTF6zF7vhB8+/Aq/J9vXfcqlp7i0OGgW5DcdRkyV3s1eUYTPMhby9UjBNQ8rl
K/Wct675AFly4yIeES8NjxG9Go789zSiRdx4rE1cp22178nI4L8cGYbpHMpgt9lV
UHnq2vL0H7jtK4JNtc+ROrSDgzprRLFfG9g9UeVfyenlbgPNq+RSRvMtr9kmLxAF
VMlfvCtD0WankUw47+yLBemtbTANIKxBECEAgAxds5qZC2txtMh+12QApjULgwYd
grWTdF3jdRUcdkCtCC07bs8WRVtn2/IHF9YjFbbHXyOtJd/J/DyObm0iepm+zzYf
KTbPCnmEfX8aBA5tvKJ21pqrp5txsnZe3SWXlHsUcdGAl5V1MHxi7PO1A+vHz7qj
HyRX6USyIx/HycDYOVFc1Oh21Cgr2V57Gt3hEq0awfwdelYDAlt848Ss1h2LANCs
Ptj7VreEFXLwwnsIL6CHu6ILi6tswHlzFdkUHwpgscgI+1JrPWdLS0qixqf5oRY8
2la9yNZT5mRD+3DuvFUE5s1p2kH2Th8jWx681P9PSWFsRUzgxtqG7+UQeXVE5BFQ
Dm27xpx47kdLgRwqGFA8ssL/s/PPDnLPLBNEFHuQYLRqRn3EslVxYKeYo299t9x7
WHN37FxrQJz+rszXP2G56nT7N8DaxzVAbYEezUoxdv3ngR4hreup+0hjciVokCi7
/vXs7W/6Skl5zWgC7K5HodLAZBAmBIVq4d/liKArndq3tcROjQN0qB8OeRy93Eh/
YwfhYuaq/0nq2Ofbww56NJ/gjP7J83T/XdUKaY1jOSG+zNZ4wTCD1iQUnBPqVrEk
Jyz6CEgsVv/wEG6lhlwVhcyfze5HJ/YSTG3pTl0dUyTC8FOrmy4D8vLX5E7cUlG/
bMNR0LsxXGxhXbSRCGMP5DmCwY7TW9FuuevuNk5VHzqc4fJTy+BpkrgvZi56Rrsf
ezkTqbOhTvSUvHMwRqa67JFvMFqApuJnl1n5OQcQRRcRDowQthnpZBZ/2UH1tn9d
cSrXscVA6sjHlzEYcNlhRz1NAfgxkHfEUtDW5aYoPw5lQPO2B9w5UyNFcmXwWIVc
UXE3Kk1rA8IlzogCcHcYEY7Fwm+Mh8WUkq7C8L8Sy970PGCp4zF+EOZ1E0dttClG
O/cBpBnyW9Zo6j5Yfgq8ibDPEY21ZJpAJN4wQtWXU/mOmL5jqVqNT9oG2J11L37Q
QBQRChEUWSpgJ6qPQRoTEeAf1OZmb9N8Q5dIqGVMoWymlIs0uetJY7x+JlBw7aLs
QjLeOS7e/O97RFEXzU7rn3B5oVURB992ZXqkOQnFkefB5HuS1L6wL1KC2mvMCEH1
xMO+TrHpP6MVc7UH6vKHny/1irYtfRyW5J1fPHKfWoGok+2Se+zTNbxNMr3Ljhzo
21y1/hEtiXUXVQn+MAktkdOiWYcOIRarMKfeERTcqzhmMBDjSakd7FuGkeemIMdg
731JOmr+X5HoECO10fh11d6jjQogt3M1ViSZfekgc14SZHaM5j37wWbkUPFOc5V8
iZ60fQhxPXR95WRVi232X+fvPaZJegthW1IV6e/HsSiOgivHY/+kHssZB2i9Ixlp
pw8o0Bnv4QZqeVPF7A6jGnwIO6Zpa9udOlrnRdytjHU/YhWJqTQJY+ZbhZHuaMds
OBE8q8BpSbc8jOKY6lPjLjyOtTRV2MHu1dAKFAyvJc1tjxiGJIDNR9CkiBdxa4Ob
jA9hLhl1dW7EHhryJBat4XV+Mp7PdKp/RoFfa7czRwtyC5548Ryjyq+NaEQRK9J1
itAOt7XSO+wOITL7nLyPGfraiZd8vEkgtfNmKUIC83/bk17csLeRxopTB0YmQ4rO
hduMlqZHCL+40mqla/F8incH4eNcH6QxNCAHPtI+fXmpUEAwIecZB/S4xPgy8teN
cVQ/Z9v7kDpKUvGuC9aj1pmBWNsXYvJB2U/IDTy2WaW6YKYnxoLwTI0Lo0fzSqSV
2E4f5WcQmZFAy1Llq2HMMmMsXRGgBk/lBluulHtMvD3eN4gKBHLLmHd7qWGvM9zr
rHu3ZGL8Mw6kGE4pOfh3pgaCV/oQgNR8AYz4bKeLq9MB7oEDEICgl2TQtFPSlBEw
EO0UUekfDdPe4lrdr7MOs0E4GZY/YQ4wFFbkHvRYhItmv34XB4CG84nJL5QLDZA0
ygNcgdEhophy4OWn6+tLVkqHWhq95KB92jjiDEYKk0jKZHOHXUBjM3BmHpRwXELk
6cDeIklnkeWJGyD4obufXiaW5mwJlBXCgv2hLF7CvEKCjaF9TDoa4Ui1L0I/R/IY
9ZGVUQeQN1CNNcc62XD8UEMdhLd+VwRpF5J7+G0aFuDaSytpKTRV/e9yQaBu9GGo
dUCwWltRTnA8AOeiihL24mzMfjx78lFmY/j3epTclCPTFUH5t8QwVYn75cP+xv/q
URJUVm3t8tH/ABHJR4ipAeul+8oVgQiRYqaMKHq3B+RKhSHFf/MTq0PUv4zbFh7M
tOxjXXKSGwFrNJyHBe6JzHRBFmXpb3StYJbYNwn0SRqMEKymC04wfZp7PJaXbthF
dFttpTZVMmkqeLC7sCC86nEQEnNWCX5HbZe1u3lfzKpS9QZk95cU0WAUeuTVrm+o
fGaPH9LWa+Hyo0OWVd1uuDMnJoLbb9DSaosD3rgHFY+DnALAUpa22RU2M5+0p0tH
b51GdziMqmbAIZr8OMYb2zWtkKLhr9fRIDqHNfOE1heVspMjvWs85Sc6vgmtwvgQ
pmfC35LspHy5tegIEvjyTwut9/i7ebEFLzplSa0vCsBfRssfnkGuooT5jAUdIGY8
5Of2hVhOzLYcy5LhqHq3nK2vFB1oXFzHN3rvqtInBHJqFlTBjVM36pKD67Prgiav
JNCyBXjVFdhbtJ/kcOovYp4h0QetRDB1oQMajMDF8MrOk8AV3028IFU3/U6SBYX0
9fEZwQGdZ6uxovoDgeCmr6CrZI7SKhdW0JufCvN3Hm2y/QZ8oMVdBcoMncdtVmWJ
VkYivOn7LvDv829WOYUhGmkS5EEX5larTlEF7q7ndAhZtuXlxIYyiB1H3JsWN9LQ
2H8pnLe48iwLqrLS1FMwhFt4Tav/wHqXoMIDGiPiujvxKdcPWDj2SPTErFwFofWk
CWGISJjIV6f9MhzXv7EwFOuv3Dbypoeufd6C8oxI1scBWMxktyiOuPEUxujZqbpl
VSgUwdn/H8NVK6WIZGdATF9Dm/7cErGwYljHCos1owZYdy3nHIaaFm/wzGs+MYfF
o83aJbe2Hg0zguplbxMF9F9L6C3u71cqAM+vPA15wAXI1AstQHUr5Rw/zGTmA9an
TDlVE0FoqKLAHow58GY2B9qQ76kQIUBJFHykPovDO6DNAl3AO8LjSO7H82ZH9W+6
aQYD22BAMCL6LEUj9l7XqX9mbY8hmn+RFYorpenuuqG1gDgwcRH7DTwAED6/YcBc
VXEiq+f0sI07s3N10CRZof6YYWtVd7RmdMJ0GG2piltJPM6zfNmwYmcbgdESYWO8
WlT5sIQiowob8bq6wZmqfEE3LwIlMagUVwWLWfs+cw/TS7ugZMdM+5Tx8akeMzva
LA6Q+MsRR2PGJH2wSuaY+BkVkYLymmFYrKhS0GfZX8K9VzOBsaS/MoW2DwYdgbGU
f5ISCzkdkLsv02x0kxGJDSDXYDyclJ3qm4zXdgwsPXD+XujlAdk8GYQE1St/LVr/
Fma10SQcalLYAQA0vESdMA==
`protect end_protected