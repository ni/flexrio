-------------------------------------------------------------------------------
--
-- File: CmacCore.vhd
-- Author: National Instruments
-- Original Project: PXIe-7903 HSS
-- Date: 02 June 2022
--
-------------------------------------------------------------------------------
-- Copyright (c) 2025 National Instruments Corporation
-- 
-- All rights reserved.
-------------------------------------------------------------------------------
--
-- Purpose:
--   This module instantiates all the logic to implement one 100GbE core
--
-------------------------------------------------------------------------------
--
-- githubvisible=true
--

library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

library work;
  use work.PkgFlexRioTargetConfig.all;

library unisim;
  use unisim.vcomponents.all;

entity CmacCore is
  port (
    ------------------------------
    -- Reset                    --
    ------------------------------
    aResetSl : in  std_logic;

    ------------------------------
    -- MGT Socket Interface     --
    ------------------------------
    MgtRefClk_p : in  std_logic;
    MgtRefClk_n : in  std_logic;
    MgtPortRx_p : in  std_logic_vector(3 downto 0);
    MgtPortRx_n : in  std_logic_vector(3 downto 0);
    MgtPortTx_p : out std_logic_vector(3 downto 0);
    MgtPortTx_n : out std_logic_vector(3 downto 0);
    --vhook_nodgv MgtPort*

    --------------------------------- Clocks -----------------------------------
    AxiClk     : in  std_logic;
    -- 80MHz Clock
    SysClk        : in  std_logic;
    -- 322.26666 Mhz clock generated by 100G Phy from RefClock
    UserClk       : out std_logic;

    --------------------------------- Status -----------------------------------
    xCoreReady : out std_logic;

    ------------------------ AXI Stream TX Interface ------------------------
    -- The following signals are REQUIRED to be in the UserClk domain:
    uTxTData0     : in  std_logic_vector(63 downto 0);
    uTxTData1     : in  std_logic_vector(63 downto 0);
    uTxTData2     : in  std_logic_vector(63 downto 0);
    uTxTData3     : in  std_logic_vector(63 downto 0);
    uTxTData4     : in  std_logic_vector(63 downto 0);
    uTxTData5     : in  std_logic_vector(63 downto 0);
    uTxTData6     : in  std_logic_vector(63 downto 0);
    uTxTData7     : in  std_logic_vector(63 downto 0);
    uTxTKeep      : in  std_logic_vector(63 downto 0);
    uTxTLast      : in  std_logic;
    uTxTUser      : in  std_logic;
    uTxTValid     : in  std_logic;
    uTxTReady     : out std_logic;

    ------------------------ AXI Stream RX Interface ------------------------
    -- The following signals are REQUIRED to be in the UserClk domain:
    uRxTData0     : out std_logic_vector(63 downto 0);
    uRxTData1     : out std_logic_vector(63 downto 0);
    uRxTData2     : out std_logic_vector(63 downto 0);
    uRxTData3     : out std_logic_vector(63 downto 0);
    uRxTData4     : out std_logic_vector(63 downto 0);
    uRxTData5     : out std_logic_vector(63 downto 0);
    uRxTData6     : out std_logic_vector(63 downto 0);
    uRxTData7     : out std_logic_vector(63 downto 0);
    uRxTKeep      : out std_logic_vector(63 downto 0);
    uRxTUser      : out std_logic; -- 1 indicates a bad packet
    uRxTLast      : out std_logic;
    uRxTValid     : out std_logic;
    -- There is no RxTReady signal support by the Ethernet100G IP. Received data has to
    -- be read immediately or it is lost.

    -------------------------------- Control --------------------------------
    aRxPolarity : in  std_logic_vector(3 downto 0);
    aTxPolarity : in  std_logic_vector(3 downto 0);

    ------------------------------- IEEE 1588 -------------------------------
    uCtlRxSystemtimerinHigh         : in  std_logic_vector(15 downto 0);
    uCtlRxSystemtimerinLow          : in  std_logic_vector(63 downto 0);
    uCtlTxSystemtimerinHigh         : in  std_logic_vector(15 downto 0);
    uCtlTxSystemtimerinLow          : in  std_logic_vector(63 downto 0);
    uRxLaneAlignerFill0             : out std_logic_vector(6 downto 0);
    uRxLaneAlignerFill1             : out std_logic_vector(6 downto 0);
    uRxLaneAlignerFill10            : out std_logic_vector(6 downto 0);
    uRxLaneAlignerFill11            : out std_logic_vector(6 downto 0);
    uRxLaneAlignerFill12            : out std_logic_vector(6 downto 0);
    uRxLaneAlignerFill13            : out std_logic_vector(6 downto 0);
    uRxLaneAlignerFill14            : out std_logic_vector(6 downto 0);
    uRxLaneAlignerFill15            : out std_logic_vector(6 downto 0);
    uRxLaneAlignerFill16            : out std_logic_vector(6 downto 0);
    uRxLaneAlignerFill17            : out std_logic_vector(6 downto 0);
    uRxLaneAlignerFill18            : out std_logic_vector(6 downto 0);
    uRxLaneAlignerFill19            : out std_logic_vector(6 downto 0);
    uRxLaneAlignerFill2             : out std_logic_vector(6 downto 0);
    uRxLaneAlignerFill3             : out std_logic_vector(6 downto 0);
    uRxLaneAlignerFill4             : out std_logic_vector(6 downto 0);
    uRxLaneAlignerFill5             : out std_logic_vector(6 downto 0);
    uRxLaneAlignerFill6             : out std_logic_vector(6 downto 0);
    uRxLaneAlignerFill7             : out std_logic_vector(6 downto 0);
    uRxLaneAlignerFill8             : out std_logic_vector(6 downto 0);
    uRxLaneAlignerFill9             : out std_logic_vector(6 downto 0);
    uRxPtpPcslaneOut                : out std_logic_vector(4 downto 0);
    uRxPtpTstampOutHigh             : out std_logic_vector(15 downto 0);
    uRxPtpTstampOutLow              : out std_logic_vector(63 downto 0);
    uStatTxPtpFifoReadError         : out std_logic;
    uStatTxPtpFifoWriteError        : out std_logic;
    uTxPtp1588opIn                  : in  std_logic_vector(1 downto 0);
    uTxPtpPcslaneOut                : out std_logic_vector(4 downto 0);
    uTxPtpTagFieldIn                : in  std_logic_vector(15 downto 0);
    uTxPtpTstampOutHigh             : out std_logic_vector(15 downto 0);
    uTxPtpTstampOutLow              : out std_logic_vector(63 downto 0);
    uTxPtpTstampTagOut              : out std_logic_vector(15 downto 0);
    uTxPtpTstampValidOut            : out std_logic;

    -------------------------------- Status ---------------------------------
    uStatRxRsfecAmLock0             : out std_logic;
    uStatRxRsfecAmLock1             : out std_logic;
    uStatRxRsfecAmLock2             : out std_logic;
    uStatRxRsfecAmLock3             : out std_logic;
    uStatRxRsfecCorrectedCwInc      : out std_logic;
    uStatRxRsfecCwInc               : out std_logic;
    uStatRxRsfecErrCount0Inc        : out std_logic_vector(2 downto 0);
    uStatRxRsfecErrCount1Inc        : out std_logic_vector(2 downto 0);
    uStatRxRsfecErrCount2Inc        : out std_logic_vector(2 downto 0);
    uStatRxRsfecErrCount3Inc        : out std_logic_vector(2 downto 0);
    uStatRxRsfecHiSer               : out std_logic;
    uStatRxRsfecLaneAlignmentStatus : out std_logic;
    uStatRxRsfecLaneFill0           : out std_logic_vector(13 downto 0);
    uStatRxRsfecLaneFill1           : out std_logic_vector(13 downto 0);
    uStatRxRsfecLaneFill2           : out std_logic_vector(13 downto 0);
    uStatRxRsfecLaneFill3           : out std_logic_vector(13 downto 0);
    uStatRxRsfecLaneMapping         : out std_logic_vector(7 downto 0);
    uStatRxRsfecUncorrectedCwInc    : out std_logic;

    ----------------------------- Flow Control ------------------------------
    uCtlRxPauseEnable        : in  std_logic_vector(8 downto 0);
    uCtlRxEnableGcp          : in  std_logic;
    uCtlRxCheckMcastGcp      : in  std_logic;
    uCtlRxCheckUcastGcp      : in  std_logic;
    uCtlRxCheckSaGcp         : in  std_logic;
    uCtlRxCheckEtypeGcp      : in  std_logic;
    uCtlRxCheckOpcodeGcp     : in  std_logic;
    uCtlRxEnablePcp          : in  std_logic;
    uCtlRxCheckMcastPcp      : in  std_logic;
    uCtlRxCheckUcastPcp      : in  std_logic;
    uCtlRxCheckSaPcp         : in  std_logic;
    uCtlRxCheckEtypePcp      : in  std_logic;
    uCtlRxCheckOpcodePcp     : in  std_logic;
    uCtlRxEnableGpp          : in  std_logic;
    uCtlRxCheckMcastGpp      : in  std_logic;
    uCtlRxCheckUcastGpp      : in  std_logic;
    uCtlRxCheckSaGpp         : in  std_logic;
    uCtlRxCheckEtypeGpp      : in  std_logic;
    uCtlRxCheckOpcodeGpp     : in  std_logic;
    uCtlRxEnablePpp          : in  std_logic;
    uCtlRxCheckMcastPpp      : in  std_logic;
    uCtlRxCheckUcastPpp      : in  std_logic;
    uCtlRxCheckSaPpp         : in  std_logic;
    uCtlRxCheckEtypePpp      : in  std_logic;
    uCtlRxCheckOpcodePpp     : in  std_logic;
    uStatRxPauseReq          : out std_logic_vector(8 downto 0);
    uCtlRxPauseAck           : in  std_logic_vector(8 downto 0);
    uStatRxPauseValid        : out std_logic_vector(8 downto 0);
    uStatRxPauseQanta0       : out std_logic_vector(15 downto 0);
    uStatRxPauseQanta1       : out std_logic_vector(15 downto 0);
    uStatRxPauseQanta2       : out std_logic_vector(15 downto 0);
    uStatRxPauseQanta3       : out std_logic_vector(15 downto 0);
    uStatRxPauseQanta4       : out std_logic_vector(15 downto 0);
    uStatRxPauseQanta5       : out std_logic_vector(15 downto 0);
    uStatRxPauseQanta6       : out std_logic_vector(15 downto 0);
    uStatRxPauseQanta7       : out std_logic_vector(15 downto 0);
    uStatRxPauseQanta8       : out std_logic_vector(15 downto 0);

    uCtlTxPauseEnable        : in  std_logic_vector(8 downto 0);
    uCtlTxPauseReq           : in  std_logic_vector(8 downto 0);
    uCtlTxPauseQuanta0       : in  std_logic_vector(15 downto 0);
    uCtlTxPauseQuanta1       : in  std_logic_vector(15 downto 0);
    uCtlTxPauseQuanta2       : in  std_logic_vector(15 downto 0);
    uCtlTxPauseQuanta3       : in  std_logic_vector(15 downto 0);
    uCtlTxPauseQuanta4       : in  std_logic_vector(15 downto 0);
    uCtlTxPauseQuanta5       : in  std_logic_vector(15 downto 0);
    uCtlTxPauseQuanta6       : in  std_logic_vector(15 downto 0);
    uCtlTxPauseQuanta7       : in  std_logic_vector(15 downto 0);
    uCtlTxPauseQuanta8       : in  std_logic_vector(15 downto 0);
    uCtlTxPauseRefreshTimer0 : in  std_logic_vector(15 downto 0);
    uCtlTxPauseRefreshTimer1 : in  std_logic_vector(15 downto 0);
    uCtlTxPauseRefreshTimer2 : in  std_logic_vector(15 downto 0);
    uCtlTxPauseRefreshTimer3 : in  std_logic_vector(15 downto 0);
    uCtlTxPauseRefreshTimer4 : in  std_logic_vector(15 downto 0);
    uCtlTxPauseRefreshTimer5 : in  std_logic_vector(15 downto 0);
    uCtlTxPauseRefreshTimer6 : in  std_logic_vector(15 downto 0);
    uCtlTxPauseRefreshTimer7 : in  std_logic_vector(15 downto 0);
    uCtlTxPauseRefreshTimer8 : in  std_logic_vector(15 downto 0);
    uCtlTxResendPause        : in  std_logic;
    uStatTxPauseValid        : out std_logic_vector(8 downto 0);

    ----------------------------------- DRP -----------------------------------
    DrpClk                   : in  std_logic;
    dDrpAddr                 : in  std_logic_vector(9 downto 0);
    dDrpDi                   : in  std_logic_vector(15 downto 0);
    dDrpEn                   : in  std_logic;
    dDrpDo                   : out std_logic_vector(15 downto 0);
    dDrpRdy                  : out std_logic;
    dDrpWe                   : in  std_logic;

    ---------------------------- Core Reset Status -----------------------------
    -- The following signal is REQUIRED to be in the UserClk domain:
    uUserClkResetOut  : out std_logic
  );
end CmacCore;

architecture rtl of CmacCore is

  signal UserClkLcl : std_logic;

  signal uResetDone : std_logic_vector(3 downto 0);
  type InitState_t is (Reset, WaitForRxAlign, Ready);
  signal uInitState : InitState_t;

  signal uCoreReady    : std_logic;
  signal xCoreReady_ms : std_logic;

  -- Resets
  signal uUsrReset   : std_logic;
  signal uReady      : std_logic;
  signal uUsrRxReset : std_logic;
  signal uUsrTxReset : std_logic;

  -- RX control/status
  signal aCtlRxForceResync                : std_logic;
  signal uCtlRsfecIeeeErrorIndicationMode : std_logic;
  signal uCtlRxEnable                     : std_logic;
  signal uCtlRxRsfecEnable                : std_logic;
  signal uCtlRxRsfecEnableCorrection      : std_logic;
  signal uCtlRxRsfecEnableIndication      : std_logic;
  signal uCtlRxTestPattern                : std_logic;
  signal uStatRxAligned                   : std_logic;

  -- TX control/status
  signal uCtlTxEnable      : std_logic;
  signal uCtlTxRsfecEnable : std_logic;
  signal uCtlTxSendIdle    : std_logic;
  signal uCtlTxSendLfi     : std_logic;
  signal uCtlTxSendRfi     : std_logic;
  signal uCtlTxTestPattern : std_logic;

  -- 1588
  signal uCtlRxSystemtimerin : std_logic_vector(79 downto 0);
  signal uCtlTxSystemtimerin : std_logic_vector(79 downto 0);
  signal uRxPtpTstampOut     : std_logic_vector(79 downto 0);
  signal uTxPtpTstampOut     : std_logic_vector(79 downto 0);

  -- Loopback
  signal aGtLoopbackIn : std_logic_vector(11 downto 0);
  constant kLoopbackNormalOperation : std_logic_vector(2 downto 0) := "000";

  -- Equalization
  signal aTxDiffCtrl   : std_logic_vector(19 downto 0);
  constant kTxDiffCtrl840mVpp : std_logic_vector(4 downto 0) := "10010";

  signal aTxPreCursor  : std_logic_vector(19 downto 0);
  constant kTxPreCursor1p30 : std_logic_vector(4 downto 0) := "00110";

  signal aTxPostCursor : std_logic_vector(19 downto 0);
  constant kTxPostCursor5p05 : std_logic_vector(4 downto 0) := "10010";

begin

  -----------------------------------------------------------------------------
  -- Constants
  -----------------------------------------------------------------------------

  -- Set loopback to normal operation
  aGtLoopbackIn <= kLoopbackNormalOperation & kLoopbackNormalOperation & kLoopbackNormalOperation & kLoopbackNormalOperation;
  -- Set TX equalization to 840mVpp, 1.30dB Pre-emphasis, 5.05dB Post-emphasis
  -- These settings selected by eye scan sweeps, but may be changed if needed
  aTxDiffCtrl   <= kTxDiffCtrl840mVpp & kTxDiffCtrl840mVpp & kTxDiffCtrl840mVpp & kTxDiffCtrl840mVpp;
  aTxPreCursor  <= kTxPreCursor1p30 & kTxPreCursor1p30 & kTxPreCursor1p30 & kTxPreCursor1p30;
  aTxPostCursor <= kTxPostCursor5p05 & kTxPostCursor5p05 & kTxPostCursor5p05 & kTxPostCursor5p05;

  -- Convert 80 bit wide I/O to Labview compatible sizes
  uCtlRxSystemtimerin <= uCtlRxSystemtimerinHigh & uCtlRxSystemtimerinLow;
  uCtlTxSystemtimerin <= uCtlTxSystemtimerinHigh & uCtlTxSystemtimerinLow;

  uRxPtpTstampOutHigh <= uRxPtpTstampOut(79 downto 64);
  uRxPtpTstampOutLow  <= uRxPtpTstampOut(63 downto 0);
  uTxPtpTstampOutHigh <= uTxPtpTstampOut(79 downto 64);
  uTxPtpTstampOutLow  <= uTxPtpTstampOut(63 downto 0);

  ----------------------------------------------------------------------------
  -- Ethernet100G Block Diagram
  ----------------------------------------------------------------------------
  -- use the same name for the instance as in the wrapper of the block diagram
  -- to be able to reuse the constaints
  --vhook_e CmacWrapper
  --vhook_a UserClk         UserClkLcl
  --vhook_a aGtPowerGoodOut open
  CmacWrapperx: entity work.CmacWrapper (rtl)
    port map (
      MgtRefClk_p                      => MgtRefClk_p,                       --in  std_logic
      MgtRefClk_n                      => MgtRefClk_n,                       --in  std_logic
      MgtPortRx_n                      => MgtPortRx_n,                       --in  std_logic_vector(3:0)
      MgtPortRx_p                      => MgtPortRx_p,                       --in  std_logic_vector(3:0)
      MgtPortTx_n                      => MgtPortTx_n,                       --out std_logic_vector(3:0)
      MgtPortTx_p                      => MgtPortTx_p,                       --out std_logic_vector(3:0)
      aResetSl                         => aResetSl,                          --in  std_logic
      uUsrRxReset                      => uUsrRxReset,                       --out std_logic
      uUsrTxReset                      => uUsrTxReset,                       --out std_logic
      SysClk                           => SysClk,                            --in  std_logic
      UserClk                          => UserClkLcl,                        --out std_logic
      uRxTData0                        => uRxTData0,                         --out std_logic_vector(63:0)
      uRxTData1                        => uRxTData1,                         --out std_logic_vector(63:0)
      uRxTData2                        => uRxTData2,                         --out std_logic_vector(63:0)
      uRxTData3                        => uRxTData3,                         --out std_logic_vector(63:0)
      uRxTData4                        => uRxTData4,                         --out std_logic_vector(63:0)
      uRxTData5                        => uRxTData5,                         --out std_logic_vector(63:0)
      uRxTData6                        => uRxTData6,                         --out std_logic_vector(63:0)
      uRxTData7                        => uRxTData7,                         --out std_logic_vector(63:0)
      uRxTKeep                         => uRxTKeep,                          --out std_logic_vector(63:0)
      uRxTLast                         => uRxTLast,                          --out std_logic
      uRxTUser                         => uRxTUser,                          --out std_logic
      uRxTValid                        => uRxTValid,                         --out std_logic
      uTxTData0                        => uTxTData0,                         --in  std_logic_vector(63:0)
      uTxTData1                        => uTxTData1,                         --in  std_logic_vector(63:0)
      uTxTData2                        => uTxTData2,                         --in  std_logic_vector(63:0)
      uTxTData3                        => uTxTData3,                         --in  std_logic_vector(63:0)
      uTxTData4                        => uTxTData4,                         --in  std_logic_vector(63:0)
      uTxTData5                        => uTxTData5,                         --in  std_logic_vector(63:0)
      uTxTData6                        => uTxTData6,                         --in  std_logic_vector(63:0)
      uTxTData7                        => uTxTData7,                         --in  std_logic_vector(63:0)
      uTxTKeep                         => uTxTKeep,                          --in  std_logic_vector(63:0)
      uTxTLast                         => uTxTLast,                          --in  std_logic
      uTxTUser                         => uTxTUser,                          --in  std_logic
      uTxTReady                        => uTxTReady,                         --out std_logic
      uTxTValid                        => uTxTValid,                         --in  std_logic
      aRxPolarity                      => aRxPolarity,                       --in  std_logic_vector(3:0)
      uStatRxAligned                   => uStatRxAligned,                    --out std_logic
      uCtlRxEnable                     => uCtlRxEnable,                      --in  std_logic
      aCtlRxForceResync                => aCtlRxForceResync,                 --in  std_logic
      uCtlRxTestPattern                => uCtlRxTestPattern,                 --in  std_logic
      aTxDiffCtrl                      => aTxDiffCtrl,                       --in  std_logic_vector(19:0)
      aTxPolarity                      => aTxPolarity,                       --in  std_logic_vector(3:0)
      aTxPostCursor                    => aTxPostCursor,                     --in  std_logic_vector(19:0)
      aTxPreCursor                     => aTxPreCursor,                      --in  std_logic_vector(19:0)
      uCtlTxEnable                     => uCtlTxEnable,                      --in  std_logic
      uCtlTxTestPattern                => uCtlTxTestPattern,                 --in  std_logic
      uCtlTxSendIdle                   => uCtlTxSendIdle,                    --in  std_logic
      uCtlTxSendLfi                    => uCtlTxSendLfi,                     --in  std_logic
      uCtlTxSendRfi                    => uCtlTxSendRfi,                     --in  std_logic
      uCtlRsfecIeeeErrorIndicationMode => uCtlRsfecIeeeErrorIndicationMode,  --in  std_logic
      uCtlRxRsfecEnable                => uCtlRxRsfecEnable,                 --in  std_logic
      uCtlRxRsfecEnableCorrection      => uCtlRxRsfecEnableCorrection,       --in  std_logic
      uCtlRxRsfecEnableIndication      => uCtlRxRsfecEnableIndication,       --in  std_logic
      uCtlTxRsfecEnable                => uCtlTxRsfecEnable,                 --in  std_logic
      uStatRxRsfecAmLock0              => uStatRxRsfecAmLock0,               --out std_logic
      uStatRxRsfecAmLock1              => uStatRxRsfecAmLock1,               --out std_logic
      uStatRxRsfecAmLock2              => uStatRxRsfecAmLock2,               --out std_logic
      uStatRxRsfecAmLock3              => uStatRxRsfecAmLock3,               --out std_logic
      uStatRxRsfecCorrectedCwInc       => uStatRxRsfecCorrectedCwInc,        --out std_logic
      uStatRxRsfecCwInc                => uStatRxRsfecCwInc,                 --out std_logic
      uStatRxRsfecErrCount0Inc         => uStatRxRsfecErrCount0Inc,          --out std_logic_vector(2:0)
      uStatRxRsfecErrCount1Inc         => uStatRxRsfecErrCount1Inc,          --out std_logic_vector(2:0)
      uStatRxRsfecErrCount2Inc         => uStatRxRsfecErrCount2Inc,          --out std_logic_vector(2:0)
      uStatRxRsfecErrCount3Inc         => uStatRxRsfecErrCount3Inc,          --out std_logic_vector(2:0)
      uStatRxRsfecHiSer                => uStatRxRsfecHiSer,                 --out std_logic
      uStatRxRsfecLaneAlignmentStatus  => uStatRxRsfecLaneAlignmentStatus,   --out std_logic
      uStatRxRsfecLaneFill0            => uStatRxRsfecLaneFill0,             --out std_logic_vector(13:0)
      uStatRxRsfecLaneFill1            => uStatRxRsfecLaneFill1,             --out std_logic_vector(13:0)
      uStatRxRsfecLaneFill2            => uStatRxRsfecLaneFill2,             --out std_logic_vector(13:0)
      uStatRxRsfecLaneFill3            => uStatRxRsfecLaneFill3,             --out std_logic_vector(13:0)
      uStatRxRsfecLaneMapping          => uStatRxRsfecLaneMapping,           --out std_logic_vector(7:0)
      uStatRxRsfecUncorrectedCwInc     => uStatRxRsfecUncorrectedCwInc,      --out std_logic
      uCtlRxCheckEtypeGcp              => uCtlRxCheckEtypeGcp,               --in  std_logic
      uCtlRxCheckEtypeGpp              => uCtlRxCheckEtypeGpp,               --in  std_logic
      uCtlRxCheckEtypePcp              => uCtlRxCheckEtypePcp,               --in  std_logic
      uCtlRxCheckEtypePpp              => uCtlRxCheckEtypePpp,               --in  std_logic
      uCtlRxCheckMcastGcp              => uCtlRxCheckMcastGcp,               --in  std_logic
      uCtlRxCheckMcastGpp              => uCtlRxCheckMcastGpp,               --in  std_logic
      uCtlRxCheckMcastPcp              => uCtlRxCheckMcastPcp,               --in  std_logic
      uCtlRxCheckMcastPpp              => uCtlRxCheckMcastPpp,               --in  std_logic
      uCtlRxCheckOpcodeGcp             => uCtlRxCheckOpcodeGcp,              --in  std_logic
      uCtlRxCheckOpcodeGpp             => uCtlRxCheckOpcodeGpp,              --in  std_logic
      uCtlRxCheckOpcodePcp             => uCtlRxCheckOpcodePcp,              --in  std_logic
      uCtlRxCheckOpcodePpp             => uCtlRxCheckOpcodePpp,              --in  std_logic
      uCtlRxCheckSaGcp                 => uCtlRxCheckSaGcp,                  --in  std_logic
      uCtlRxCheckSaGpp                 => uCtlRxCheckSaGpp,                  --in  std_logic
      uCtlRxCheckSaPcp                 => uCtlRxCheckSaPcp,                  --in  std_logic
      uCtlRxCheckSaPpp                 => uCtlRxCheckSaPpp,                  --in  std_logic
      uCtlRxCheckUcastGcp              => uCtlRxCheckUcastGcp,               --in  std_logic
      uCtlRxCheckUcastGpp              => uCtlRxCheckUcastGpp,               --in  std_logic
      uCtlRxCheckUcastPcp              => uCtlRxCheckUcastPcp,               --in  std_logic
      uCtlRxCheckUcastPpp              => uCtlRxCheckUcastPpp,               --in  std_logic
      uCtlRxEnableGcp                  => uCtlRxEnableGcp,                   --in  std_logic
      uCtlRxEnableGpp                  => uCtlRxEnableGpp,                   --in  std_logic
      uCtlRxEnablePcp                  => uCtlRxEnablePcp,                   --in  std_logic
      uCtlRxEnablePpp                  => uCtlRxEnablePpp,                   --in  std_logic
      uCtlRxPauseAck                   => uCtlRxPauseAck,                    --in  std_logic_vector(8:0)
      uCtlRxPauseEnable                => uCtlRxPauseEnable,                 --in  std_logic_vector(8:0)
      uCtlTxPauseEnable                => uCtlTxPauseEnable,                 --in  std_logic_vector(8:0)
      uCtlTxPauseQuanta0               => uCtlTxPauseQuanta0,                --in  std_logic_vector(15:0)
      uCtlTxPauseQuanta1               => uCtlTxPauseQuanta1,                --in  std_logic_vector(15:0)
      uCtlTxPauseQuanta2               => uCtlTxPauseQuanta2,                --in  std_logic_vector(15:0)
      uCtlTxPauseQuanta3               => uCtlTxPauseQuanta3,                --in  std_logic_vector(15:0)
      uCtlTxPauseQuanta4               => uCtlTxPauseQuanta4,                --in  std_logic_vector(15:0)
      uCtlTxPauseQuanta5               => uCtlTxPauseQuanta5,                --in  std_logic_vector(15:0)
      uCtlTxPauseQuanta6               => uCtlTxPauseQuanta6,                --in  std_logic_vector(15:0)
      uCtlTxPauseQuanta7               => uCtlTxPauseQuanta7,                --in  std_logic_vector(15:0)
      uCtlTxPauseQuanta8               => uCtlTxPauseQuanta8,                --in  std_logic_vector(15:0)
      uCtlTxPauseRefreshTimer0         => uCtlTxPauseRefreshTimer0,          --in  std_logic_vector(15:0)
      uCtlTxPauseRefreshTimer1         => uCtlTxPauseRefreshTimer1,          --in  std_logic_vector(15:0)
      uCtlTxPauseRefreshTimer2         => uCtlTxPauseRefreshTimer2,          --in  std_logic_vector(15:0)
      uCtlTxPauseRefreshTimer3         => uCtlTxPauseRefreshTimer3,          --in  std_logic_vector(15:0)
      uCtlTxPauseRefreshTimer4         => uCtlTxPauseRefreshTimer4,          --in  std_logic_vector(15:0)
      uCtlTxPauseRefreshTimer5         => uCtlTxPauseRefreshTimer5,          --in  std_logic_vector(15:0)
      uCtlTxPauseRefreshTimer6         => uCtlTxPauseRefreshTimer6,          --in  std_logic_vector(15:0)
      uCtlTxPauseRefreshTimer7         => uCtlTxPauseRefreshTimer7,          --in  std_logic_vector(15:0)
      uCtlTxPauseRefreshTimer8         => uCtlTxPauseRefreshTimer8,          --in  std_logic_vector(15:0)
      uCtlTxPauseReq                   => uCtlTxPauseReq,                    --in  std_logic_vector(8:0)
      uCtlTxResendPause                => uCtlTxResendPause,                 --in  std_logic
      uStatRxPauseQanta0               => uStatRxPauseQanta0,                --out std_logic_vector(15:0)
      uStatRxPauseQanta1               => uStatRxPauseQanta1,                --out std_logic_vector(15:0)
      uStatRxPauseQanta2               => uStatRxPauseQanta2,                --out std_logic_vector(15:0)
      uStatRxPauseQanta3               => uStatRxPauseQanta3,                --out std_logic_vector(15:0)
      uStatRxPauseQanta4               => uStatRxPauseQanta4,                --out std_logic_vector(15:0)
      uStatRxPauseQanta5               => uStatRxPauseQanta5,                --out std_logic_vector(15:0)
      uStatRxPauseQanta6               => uStatRxPauseQanta6,                --out std_logic_vector(15:0)
      uStatRxPauseQanta7               => uStatRxPauseQanta7,                --out std_logic_vector(15:0)
      uStatRxPauseQanta8               => uStatRxPauseQanta8,                --out std_logic_vector(15:0)
      uStatRxPauseReq                  => uStatRxPauseReq,                   --out std_logic_vector(8:0)
      uStatRxPauseValid                => uStatRxPauseValid,                 --out std_logic_vector(8:0)
      uStatTxPauseValid                => uStatTxPauseValid,                 --out std_logic_vector(8:0)
      uCtlRxSystemtimerin              => uCtlRxSystemtimerin,               --in  std_logic_vector(79:0)
      uCtlTxSystemtimerin              => uCtlTxSystemtimerin,               --in  std_logic_vector(79:0)
      uRxLaneAlignerFill0              => uRxLaneAlignerFill0,               --out std_logic_vector(6:0)
      uRxLaneAlignerFill1              => uRxLaneAlignerFill1,               --out std_logic_vector(6:0)
      uRxLaneAlignerFill10             => uRxLaneAlignerFill10,              --out std_logic_vector(6:0)
      uRxLaneAlignerFill11             => uRxLaneAlignerFill11,              --out std_logic_vector(6:0)
      uRxLaneAlignerFill12             => uRxLaneAlignerFill12,              --out std_logic_vector(6:0)
      uRxLaneAlignerFill13             => uRxLaneAlignerFill13,              --out std_logic_vector(6:0)
      uRxLaneAlignerFill14             => uRxLaneAlignerFill14,              --out std_logic_vector(6:0)
      uRxLaneAlignerFill15             => uRxLaneAlignerFill15,              --out std_logic_vector(6:0)
      uRxLaneAlignerFill16             => uRxLaneAlignerFill16,              --out std_logic_vector(6:0)
      uRxLaneAlignerFill17             => uRxLaneAlignerFill17,              --out std_logic_vector(6:0)
      uRxLaneAlignerFill18             => uRxLaneAlignerFill18,              --out std_logic_vector(6:0)
      uRxLaneAlignerFill19             => uRxLaneAlignerFill19,              --out std_logic_vector(6:0)
      uRxLaneAlignerFill2              => uRxLaneAlignerFill2,               --out std_logic_vector(6:0)
      uRxLaneAlignerFill3              => uRxLaneAlignerFill3,               --out std_logic_vector(6:0)
      uRxLaneAlignerFill4              => uRxLaneAlignerFill4,               --out std_logic_vector(6:0)
      uRxLaneAlignerFill5              => uRxLaneAlignerFill5,               --out std_logic_vector(6:0)
      uRxLaneAlignerFill6              => uRxLaneAlignerFill6,               --out std_logic_vector(6:0)
      uRxLaneAlignerFill7              => uRxLaneAlignerFill7,               --out std_logic_vector(6:0)
      uRxLaneAlignerFill8              => uRxLaneAlignerFill8,               --out std_logic_vector(6:0)
      uRxLaneAlignerFill9              => uRxLaneAlignerFill9,               --out std_logic_vector(6:0)
      uRxPtpPcslaneOut                 => uRxPtpPcslaneOut,                  --out std_logic_vector(4:0)
      uRxPtpTstampOut                  => uRxPtpTstampOut,                   --out std_logic_vector(79:0)
      uStatTxPtpFifoReadError          => uStatTxPtpFifoReadError,           --out std_logic
      uStatTxPtpFifoWriteError         => uStatTxPtpFifoWriteError,          --out std_logic
      uTxPtp1588opIn                   => uTxPtp1588opIn,                    --in  std_logic_vector(1:0)
      uTxPtpPcslaneOut                 => uTxPtpPcslaneOut,                  --out std_logic_vector(4:0)
      uTxPtpTagFieldIn                 => uTxPtpTagFieldIn,                  --in  std_logic_vector(15:0)
      uTxPtpTstampOut                  => uTxPtpTstampOut,                   --out std_logic_vector(79:0)
      uTxPtpTstampTagOut               => uTxPtpTstampTagOut,                --out std_logic_vector(15:0)
      uTxPtpTstampValidOut             => uTxPtpTstampValidOut,              --out std_logic
      DrpClk                           => DrpClk,                            --in  std_logic
      dDrpAddr                         => dDrpAddr,                          --in  std_logic_vector(9:0)
      dDrpDi                           => dDrpDi,                            --in  std_logic_vector(15:0)
      dDrpEn                           => dDrpEn,                            --in  std_logic
      dDrpDo                           => dDrpDo,                            --out std_logic_vector(15:0)
      dDrpRdy                          => dDrpRdy,                           --out std_logic
      dDrpWe                           => dDrpWe,                            --in  std_logic
      aGtLoopbackIn                    => aGtLoopbackIn,                     --in  std_logic_vector(11:0)
      aGtPowerGoodOut                  => open);                             --out std_logic_vector(3:0)


  uUsrReset <= uUsrTxReset or uUsrRxReset;

  -- Synchronize and delay the deasertion of ResetDone and Ready.  This mimics the behavior in the xilinx example
  process (aResetSl, UserClkLcl) is
  begin
    if aResetSl = '1' then
      uResetDone       <= (others => '0');
      uUserClkResetOut <= '1';
    elsif rising_edge(UserClkLcl) then
      if uUsrReset = '1' then
        uResetDone       <= (others => '0');
        uUserClkResetOut <= '1';
      else
        -- Delaying the synchronized reset to mimic what is done in xilnx example cmac_usplus_0_lbus_pkt_mon : rx_gt_locked_led
        uResetDone <= '1' & uResetDone(uResetDone'high downto 1);

        -- Release Reset to Labview after aUsrRxReset(probably superfulous) is done and alignment has finished
        -- Release it as synchronous to UserClk
        uUserClkResetOut <= not uReady;
      end if;
    end if;
  end process;

  -- This small statemachine goes through a basic initialization sequence taken
  -- from a Xilinx example.  The sequence is
  --  (1) Wait for clocks to come up and stabilize (uResetDone(0))
  --  (2) Turn on everything and send RFI
  --  (3) Wait for the rx allignment to complete and then transmit normal data.
  -- Note that waiting for RX Allignment takes 120 us in simulation even when
  --   SIM_SPEED_UP is defined.
  process (aResetSl, UserClkLcl) is
  begin
    if aResetSl = '1' then
      uInitState                       <= Reset;
      uReady                           <= '0';
      uCtlRxEnable                     <= '0';
      aCtlRxForceResync                <= '0';
      uCtlRxTestPattern                <= '0';
      uCtlTxEnable                     <= '0';
      uCtlTxTestPattern                <= '0';
      uCtlTxSendIdle                   <= '0';
      uCtlTxSendLfi                    <= '0';
      uCtlTxSendRfi                    <= '0';
      uCtlRsfecIeeeErrorIndicationMode <= '0';
      uCtlRxRsfecEnable                <= '0';
      uCtlRxRsfecEnableCorrection      <= '0';
      uCtlRxRsfecEnableIndication      <= '0';
      uCtlTxRsfecEnable                <= '0';
      uCoreReady                       <= '0';
    elsif rising_edge(UserClkLcl) then
      if uUsrReset = '1' or uResetDone(0) = '0' then
        uReady                           <= '0';
        uCtlRxEnable                     <= '0';
        aCtlRxForceResync                <= '0';
        uCtlRxTestPattern                <= '0';
        uCtlTxEnable                     <= '0';
        uCtlTxTestPattern                <= '0';
        uCtlTxSendIdle                   <= '0';
        uCtlTxSendLfi                    <= '0';
        uCtlTxSendRfi                    <= '0';
        uCtlRsfecIeeeErrorIndicationMode <= '0';
        uCtlRxRsfecEnable                <= '0';
        uCtlRxRsfecEnableCorrection      <= '0';
        uCtlRxRsfecEnableIndication      <= '0';
        uCtlTxRsfecEnable                <= '0';
        uInitState                       <= Reset;
        uCoreReady                       <= '0';
      else
        case uInitState is
          when Reset =>
            uCtlRxEnable                     <= '0';
            aCtlRxForceResync                <= '0';
            uCtlRxTestPattern                <= '0';
            uCtlTxEnable                     <= '0';
            uCtlTxTestPattern                <= '0';
            uCtlTxSendIdle                   <= '0';
            uCtlTxSendLfi                    <= '0';
            uCtlTxSendRfi                    <= '0';
            uCtlRsfecIeeeErrorIndicationMode <= '0';
            uCtlRxRsfecEnable                <= '0';
            uCtlRxRsfecEnableCorrection      <= '0';
            uCtlRxRsfecEnableIndication      <= '0';
            uCtlTxRsfecEnable                <= '0';
            if uResetDone(0) = '1' then
               uInitState <= WaitForRxAlign;
            end if;
            uCoreReady <= '0';
          when WaitForRxAlign =>
            uCtlRxEnable                     <= '1';
            uCtlTxEnable                     <= '0';
            uCtlTxSendRfi                    <= '1';
            uCtlRsfecIeeeErrorIndicationMode <= '1';
            uCtlRxRsfecEnable                <= '1';
            uCtlRxRsfecEnableCorrection      <= '1';
            uCtlRxRsfecEnableIndication      <= '1';
            uCtlTxRsfecEnable                <= '1';
            if uStatRxAligned = '1' then
               uInitState <= Ready;
            end if;
            uCoreReady <= '0';
          when Ready =>
            uCtlTxEnable  <= '1';
            uCtlTxSendRfi <= '0';
            uReady        <= '1';
            uCoreReady    <= '1';
            if uStatRxAligned = '0' then
               uInitState <= Reset;
            end if;
        end case;
      end if;
    end if;
  end process;

  process (aResetSl, AxiClk)
  begin
    if aResetSl = '1' then
      xCoreReady_ms <= '0';
      xCoreReady    <= '0';
    elsif rising_edge(AxiClk) then
      xCoreReady_ms <= uCoreReady;
      xCoreReady    <= xCoreReady_ms;
    end if;
  end process;

  UserClk <= UserClkLcl;


end rtl;
