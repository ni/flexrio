`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23616 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
FVgMhmFuxFvYsi+npZjztKZidQFVaz+CqA+G5oMIoDlz5pEyquDJQR4W7Rt/OKTi
fqFUk/+Rfd80kXCdQoF6aCpV0KqtyAcfXA3/adhZdXavXyQ/jk9vAXhcTeSzbztm
43xq5EMUzhoVBwL0ULRs2KOB44i34I3CBXqIU0rYCA7M4jVJOJcyE/JcD8cMFWva
rknQOWYWBDMoVJAJShJIVqSkrW95Sx6a8ZK5UZmeq0eLTKnQ/+5Rhp/S1Su5CF+M
08tWj+eSNQcgIcIRAkRTPeQp5/EH+Fba8RJxJ5akGIvG1b4UGEj1dyYvhlFPhnaS
rcGeRJv3RF7WCNfP8pUTi9sCnQ8sHYuQnGT4S1A9AUykHY1BK6U0eOd52Tmcvxme
Xvs2ZoQEL+pjqkWTXvrNEeY/HvkCip7vBejXkBT0ir8lVEt/QlpM2SAUTQX752+z
lfMWldkm4YfCc5LcbE57lHg1Cts0KsNWtpnfLYIKWnB0wX6ip6/iWYFW8Xpguedy
TF0be0KO1Qb3MZuP1gDH9F65oGDnOLYpEQRX+hqyhzjHdlaE9XRZTKQ/Czb7WB94
r56XVdiYFFqDfTNd1cV/h3b+3BPb0R15rqkJSk/HTfyVNVvnrIpFmBp1JOa8W/F4
F4hnMgKCTT1tOsX26/NSIGccGnna98F6/mI96czbnYW+AvlmyoS2I+9EdGUNNYIC
ZpdWj6j3rupzq/5SaZXXZ9FSBEifU97QDiRR5tePa+Ktt10+N6W+R2I9/T7wc93w
LJCWsA46vdQtpZFF0W3V+1Ho3cGCAYbmSAzoDpMrKJwP4vMdI7b5O8Bo/o1xzQN4
u8tmWKKoNR+1q3AWiBv+kHniU9Ychcy8QdEW2ccnzg1J0LzhPqE6QTG2L8MBvUKh
E0kPcZNLL8nFJCNRsNB4rFmQWBVTL0gP3fsGppS7yeFWJI1cw9sODCoHJVizzAkh
6QFsLRnnajMgq/tcxpltFS5KQheb6up5x7EyG3eQQU9eJX/0ryEWvkJyO4q+NSSY
E1hbE6iYFCW6imBewOA1ctwWTWYz0WGtcnph9LSF/wYsLblQJAG+iIyqwK6lhhB/
DjTCOMngrsotF/T9VJ7gAlKWnnGF4vaBEk7XXortOZmsUaKHmlc281FugrSZuYwA
JsN84vMa/SVQEkBsch7vXW1gOhy3UGVnACK5TLPAlG+qR5oBXdiBa4ML3uZd+ReQ
WinIsG0nCO/Vbw7pU1AT9Ut92Q8QPIi8B37T2uMhEHFbvXH+2k+SqrWL0izOKiZc
/9iX0FvO9IaCpufLvd3zFXFEsp3hc10ix0n3na650Ln/tPLJvJ0xmOC58FbEeoZD
m+8oZYa3S3xVdf/xv7crvsiQfoNWJkPWY8Cv4ppcvVCbyC2MBiiqQkRZv8rur0ht
e25FJiVbAUYwilZ5izQzbEt+5K031iOWNrsU1pkrhX7HHYuF2lvF6SMsyMG6Ptbc
cF0bppCFxnJ7nwUvGwtXqAIDJhA9AeJ4AwyuyuFCTGYk0BtMVZRsAqU2GaXqQBen
ixrItvd0WqG4yDiS0JHpWQX/rerFqWLgR3VtLxQ66IKEAZxktO0UCeg41AuypmNz
FuV/tW7Qa6WDBHFW3EW160oEN2BhgOR3c/Vg+5yqqdnPaZwfudMRbWZ65iN/FgTi
Lm2ZwLohCKwWrUTJ/8P44uUK5ccw/Xliie+5Un6JPtIvOEELHdf8J8MU1N5dCmsc
c/cjFARRb+tuQHpxUi2LSGNIXaw7L2z+yiGZ1oqgNcmpLmFD8Tk5Wdb+f4frEdog
K1VK+xcoMfOwxCKTla7/9no4wJ5i6r0Ur7ExEOAc5eOUo9y3SMh0boGTBIIAuF+3
PS2cpy4YxMr9E9ZoQAhn7fAVyeF/ykOJhxPan3cFel1T3FwNYS54jniY3IhP77M0
qb+OdxiPwUBO1qox5gPQsWTtndQVDEhTUqEdg2ad51vIDCRKW6t194yEVqq7guBP
jx0qGVwB8iwZB1KhqUdNIoGVC4hfJWFYbMaf5qGAsx53umMXvSpCjuVv1CnDmDnP
zMynox8qd5Ml4CTK4q4624v3yZeKC6Np+mnmF6XR7rcRHQxv1IJZfBKuYVA6ccYy
EU7PEzmfPr/dxOOT3/RY01EMna6zuLqF5CO5W13PPIcZ3EvSq6gGexLDj3vpajDm
BY7OsvwumSSiafEfg+xpuqSsdG9M4hroRNCwqdERqlksSO+leMHNAXDW0F5yQQTc
oshkH7Mi8ztFdpgiqUepkacsOxdLWCUomPo50DyDj/1fhd3KQMYYjvee6pSSjqJ9
Vew0rwdPgWFhZOPEpRc0k865GcqPE+ItHwRYXFRVZV9Xij/AAZCt5h9YgZczxHHP
8AKmrKB+k57d4YkUJmWC/VVy6vC4AnN4tADW1tnyzRrz1cdtGFY3pzy9ep1ZnJ3W
5bCdbkutgwoP4TTsC+nB9T3gxjTG3IOWi+t630xI2z0GUh8Arf3OWbMdh7cVC/o/
b3Cb7EbFuQoTiIrvAa+xj0DKnjPwWcY6EDEIPKkNPQiWkDIIDJJqlycwTQ2E1nOH
xkkudhABLDwEeJzHrbCJxkBmNexhPx7+AhPQa1JWaADxiE29Dbs9WVq+n5CN9AI7
HCZ9pU3m8dpCH11gFl+vcilROICfNoK3mjS5vhzTUm4uKjq/i2yFMpD3aCmFRX6f
42JtnLCqBkkz2PuDa/xHBlMSejJ/jYwOQM62ZntSB6kKtGrKDboARQQa2/BWw/yI
ki9dZ+ywMZbsCeEBnLxmGIs1LNSO6wSbqzUDmfD7XY4PNHrdgzVzq58qozycNFtd
1852Az7cz7aeoX32N1CRM+HtXbLAKEp2/9xjXVPQKuSdyvB/Ok4sNrvkcWrZqVYW
TfnSH7zopp3oKlXsiFPL+HJjuLRNQQNtiTDoZ2IyofiT5HfNKsJL7Z881s/ojd0d
acdb4+iAHVnV8IcfjfZNihCXoTEQGgF2k4OkUCReLHO8BsweKjQHPYD3R94LAdl0
nGQILImEe+oqbgQR3/4YAOyTMbG4f+2FX+0trF6N68xLJ4yx+2jA+FIcZRxVywYp
xqsIBT0gk0If6NDF4EuW/kzTdm0fmpu/+ogTFD740cccCviDL33wCIRNGkaiD1pr
voRG9JFtcSeGVeapFqNvNv/iZM4ALkLhhzP+TGCXviota1D/n3d8InbwQvQpn0I0
QB2gdPz3ybm+HqIFBSxWbArDrT8AyXeQ69KCKEQexHkDO3R5hqShpGjQaslruP2b
MTSXbbfnx55hcPbd58OhOp16Cgnn6dGVOqMrqps73KaCXT4Uc/iPofMD2N92gSra
aQ61F6JgLCf/Dw50njIZwfpGWrryvqL6GHKAYoFrH+S+KIWNffIjJPO7MwaqNBzB
7cdmr/8OeBEPayCQ13B6Xj6bqFJ8cXoHFTQPb5EvE4grqaODjBMpZOYVgHoPrEMi
H+RqD/yWOv0h0kMDPzNjpsAAVkL46IoluBuSStTGJEFJrV/WJXQ/YIpz44dI8j1i
pS7lj5xz+0vWqQYQAjpRmaLVllWMsxB+b7PysdyhxSvruD/ATn8sTmrWX0Pg4Gzj
NkBXlXbzk80n34WxFUzVgqyxevVDOtnlUjgwkb+QKA3dFJh6i7i/to3rrRd+4cP+
63w1R94h6v6nE75JmN3vYVoSOWprFqiWeNYevKsfEYn8wFbd3SDEoH8WWM+dgzfj
Kdd1vNfjWGOTCoqzavMUgka4zQjKnY209WTk5G2roFOmmspk5e2wM1prnqKC6v02
p4ZdqiNJVvESu60EGZFNY0KCQNk7oiIzaM0+tfHwdnFkdBMa6YxCqi5VQ4zGXUwh
o9MVD3DCpDVdVKC2D+rxp9DZq1aiCMGSk7oqnoIrbeiEZjK5VL89VwuOaKW6TFW/
5/t2FIq7ImXuhsqRePpDFSiEdVz5djl+Pn8IjmFY8cuQFkMPWPTUMcasBeFeWmc/
+J4OVAy0LA1zgWITCZ4FltGTu0R0FTLeVI/yQQkEiISEN9b+2IstLA+PQ5BmRiKO
V9IxaCtmgXS/wJSlJ/ZN0DCWJMtTtoUi9qq+n/Gb8mPCWut/HPZ8m8i9Y8uIN2Mc
1sGspFSDn+CL4E901NCC3nawddj9lbf1FCwQlhv3+KnXDkB8maeaGlOs6LUG/urW
PLJxUbB5ynCOQeYbTXC6a1BCQzV/fhSn23g0FNXWBldLwSH9l8DX26Mn3Z/6+Upy
y7f59omgiyTaQd9Y8YaBvojKlDu9nlotoUNHjW66VD0tqtWZwrbaQl7ieFwCbxmi
cb9aGYsU4TFQBQIwQ2uKOIgYYGzaZWuUyDBZ4Q4jEshrsuLuR7uz78wmTwOD51cs
uZYZhfDGoACrfRkUZQKqNuGQke9H4cwBUlQjFoXn55NZJREkg9J8Q0b5PgUhRaH8
dGtsC++xpts/t8sQ45QYOlhRKwfInyTUuTSL4GcUwFWOEXNp0TcZHxA/KCxzPham
+/tnCl8tiV5ulkN7ru33e4VHOoUvlTqLTbhRL82PDZfHtAX5bA4Pl6lr6PSQmNBd
tUEgjvD1qNGAWfS9MJ08Ie0g7NlovZZi4AnALq/bAnOIF1gxFf2lvRiBnNoVtUPE
ga8lexpBAGzNQBapKFfREeWDNCBySwfr0M/gTYhAGWVEroVpTX6m9CyBWRZabuyL
aSKkZ23IJ6Y5DnlOm8K79Iw0hmYLQQaD0LBCG+ThUMbGVGzO4e1HRovjI/uhVZzy
Uzcoylq5Gglnb/zrlipS9srWoBsHe7MuNPqETk3pV/hy0cYAW2WtGDCeRgNP1e/0
Mg0cTyruMoZCsq15LlbawvAe0WvFuyDSM1Um7xQpeg0+wg0j0ITf8DJCZvQ33X11
vAqWKPET3Fy5B2SRG7UZwI9KX8YVz/xkjqIuDhzbT8uTrHLl34clfJUis9ztRjZS
lFsdWwp5zDpYKGV8Lu7TP5kqVMdE3d5LnVolIzJPY1xtj1158UEm39ziAJ+/Yasz
tgqXdLyjcTs0yy17n0vVW5vXEM6TgiZhCs9VLb7YAr4D6WEFwSkpnWxj+VwziCsJ
68ViVXr+yGswiJNoHYTJD/6/8xxYe6VDgP1M/6hRwMx5pQYrZKvuJIwdWTYG9FB1
4SzEHH/nbaTXzFOMByBF9Ku5hY7iI90rjx/7Fwf4kdJ33y7FQKxUU39IV4PziPkG
mFHhftBysbaujr78W5Vz3kgM23e3O35tFcAeM95DLi4qS+kdcUBBKFrHrqDW4fAx
xxt8Jgv1SWBuKAeS0KXBAuAotfzNsGfNkmeBP8mdvNC/ylkCRKMUgofPhr17GtbF
engCQSa5QsxE5uXOIYTc9i7OI2dgQKTgzO02ef1+Lz8IOixqkYxSybfFheE5rD2t
gu4wXlRrA8abGMVHd5TGxfOrCdpJj0xBW4pfDh55QyiAy7UaMfA8hmLEWtgfK0vK
QRyoM/2e94HF+g967w2JOP8b3zFRgqhC/bRcaEYe27Yzhgy5xhTHr81+3ruVKbrR
O/BYW7T52K7fB/mapOQ3L/5S9Se6id/KDwPMICuSq/oKfSgYcKOlhxW4IUDLwZeS
n/6f5JhFKiUXIwAy8jIqGRJdwrpUf1a0o54Fne3SSyWDTUNM653ER0YqYVr9zlXw
WpiADYGtHHr2g5OSSvgqTHn/vHMndutToYXoS5pOsyJjDdCwQ56/irFLT/7x4TtA
CWWWGgcyEx8NwbeMcQZ4RJUlL4KuHVvKjbo7ZF3nG38EuMJzKKe9dcdYfl6H+n9/
OVFa8DqONYAlxNp548F/MFJ9CGk17XOFr4rSnn52un1DxakfqE3Yxa3F2R/Ofr2E
SJDHzDH883imlpFoD1QlEgRpt0Mnkp2XuCwBwznRtmeewj5IYfFQbTLB7SDNRbfl
O+rU1OFzH/gVYA8ip2yHYdSNYtjmHViT9tbrqi2GPtj/wlglaAN144K8QRbXAIly
a2NHM19yN/p5rfs4b6TnMNx5nLO71Wa49cdcHQPk2xDWWHxJndqfC2WBHKqVGjrl
/vGlNuTZcEITI+QyABc6A94/AOslx5ZFeAEywSMFfs6u/yKdmcB/fsVl3g3hT9lZ
SryA/mX8EzIh8WV0TzEeacXnJtwj4wg95yby/YEXfmWXZjGSRZ3IGbXWSXL5viAd
p0Vw22CDyi7q1Np8V0Lo0Ll6/puN9FeCu2K90oLTMjy+P1lNOpmfCEz7G9dUCAjz
2WwdWtyEC8bURBZRVCJxIbJ6K6etVxAkecLTvdkTeXgmuEmbGS2eInKGXDHxZTJF
/e+kK+FDT0OsrommaakaQue+zVlfnscNHVlDktdLSkFYiQ8ebjdZRPbCQrAvLQQ5
b0+NLVN7Q0yzoB87Xd4/xUxkQJeqlsj739LX6RbRzSZYn3QXi0xVQIGfpuKgGs/m
T89jzPk+FINfqD/XGzEf0sLEEU9tQBWBoc0BmxwCc4T2Og3yB2uTXE+Fop6gSgf/
04l0PiE4JQ3Hl9dsi8buaBew0Pfz9o6c0E5+mcOYgMvMN7asm038vOZt0nghz7uG
Cpn4u4f5M+Ojczrgsns8gWkODuiJ2lVhp3IU9JllkVzTOdYGeKnRsWcHtTM8quGO
g+Y0E2gMZM1BRTIdwB4XkjUVKn1TK6BVFvFX1iiNJoXlndL8NNw9zTytUh/Qgc36
t/6lPyIcGc/o4G+UgH/sAeJI+qxinj/MSyJhsYvL6ooGDH0CrWf25nDLHEB3iMYx
8wKR1mbCGY3IPlsNS9lwt4UOpaD92IIj0epYlZ7mtw+8BKTjhIcQrCrXXcbqvQ8M
mKeqXbwLDDtnCBH5fXLD3Qyx2WORtvDxzNT2zyQnYS0GtUr9GlJAdDdWtZJ2Cfft
StymDYBBkNFHV45i+QB7M3YNyI8jQpHQWTJL/C5+wddlg2p82CZbRESN83GYlz+S
bKpAyAKpYWN4EVeyw8b1PYIWoJqNaAms1d9oDiizY0sEH+tNq3/s9tyXZEgVg6ME
dAQu6vC2/O1PR6o4MzTG9J97Wfa8dmTa92N3K+6W9ghQ8Qjfpj48vwqqtiNQL1KZ
49ZNC5+YXo2ZdhYtJSz35neH4gtKArhoqVgEDiFqhNExS77uxaX2gAHUa6Vts1JF
7BCd2pIC/JlzCrRNwyRFDmMSzPvuFAIIQGW6xvXF2DzHRKE4k92DY7UmYFmFX1yY
/1NhFwpRpQMiGVLBpWhwWtCV37FMSY+t1EIxN5jsEs4PP2vylbKNL7xrEoqSTFCZ
h97a2yKLsPmg+mPecUCGbOqymqpxQz8vP1HEz9RB2j1rivfJbLRZVd90r1aoYT+i
uN0cCXzJgM1/NZQfALTVmoeV07sdbCo6qI06lB+Odb+XXTeOap0qHCzCOyx9zav/
/9al1Oe8d7xRAELKH4q06kJMwpTSoQV84BN4Bvhrf/nKj1i9dzlslUI00EWz53mx
r2YFhRn5vX8HYCbuFlb/jn9U8pJwej0LM9SmCr53LA0Pwrsd7shZKHxWFgeDdfSD
xoWFUmycAPwr2oIqem+Jay/WWKMVGl6n/8phAgb1QIriuK4RG16m7S3Xj33FFdYp
NpwP1bs3VaXYB2zZznCEDG4gdfgGdIXs14I+MIeaYZJ4Mpphnw+jrh8Gk+4KKPFl
EhBVQe6c6CriqHZMnQUqE6NCdMEKqlS130xv2rmaKNWC+j7KHFIbMVex8Kc4VZW1
4MoTY+3i1xxAuwEn10z5yqt/SiaOK3wzGDDcwaMU91gnGw2y+/NB8E0FSwnh66Gj
7hhRk0bcdBBKQmzj2eOZ2MYGTZ+K5LkjFaJ8AkJ0M7ovyfYHZIsQlAWBLz0Vul3W
vctE+wfcvBcWE4deE4lRssSVul2RBgleZ+dfm+swgvaCMT2FgF01Rwv9i3BUfooO
43xrRop6WR2BrAEykK5wXEPGq6emQeG3XyXYHpTPJloxyrycOP4Qw9OJNYUGTjcF
FWjH0KjYkIJ+wZl8MUbjhdiJI4PTW36XLxtr092IitGEDs3cowrxYYliRRwMdKXi
TMbHr7jODC+OEod+lajtU40BrN0FiOii503aM8gVt/OIMnQ55XMF+2+jna02LZpN
J20hLktQ6BtsKAQDNOWRsa3CXU7by+/Xt3MnT8qleCsjqtknAr6EsqDGKzYE+KLE
WGpGQ0EUDY4FBvH3R6OwcU4iRu/FMnc4dMTHfWE90m1kC/ufY3Uq3QjUVrs2U6Kc
RQoiSfB7vhW5pLRRP2KNJvqomBuhSaCErsNvNTKUhT/UfIoL2KcSEYM0aJXR031U
1JFYo9f3+IPRe+Hu+lqACoy1FFCER44/iaFQbLSr4p3Gl9M1Pof3emnYusPwK4KT
CTEdr9YiL2x1+zaC2hgC95zUeTRcJCNQZL73FIh71J41siGZwYihLYDRirDUFuAd
omVBLLikdOtaG8BYzJN6vehWArH4dy5JCBNP1+T3uWfn/HKUZZ3EfdM+FOwBQqcj
sz/O6L4DHYCjHhpdQjpOm/4i9s3fBea5cnIzneVXUlolOot7NcmRfzrg8FIkev0/
sn+OY4WNS7GkNrs0LNkFBxJJLv+srVsbvgQPZCZpYcG5y2jJOhbFx4/oMeY5Getu
ALuAavI9svZ4Dox9pSGePXJroB3FyxIedaHdboS4D0JcFjDAzMvY4gF7AeDwy+JS
1lKoLVj6vItKEZNEd1Uv5aHFdFlOd277aEE5hmReTeIzY3t0/Afg3ZtQotmi+Wfa
5hChh6z0CJMNAfavNV/tpu99UQ56nNa5fMFgpdLtSsu9JILJfvE7ZAb29gfCEwbA
KDrvswSekuouTf5R1nBKc7M+kROtoZk0KLK5YAh+31wlj7VGT6uMshe4vpbZ+mLV
DQ4KwtIUySunoXwALC+otXfybuvjLQ4QDQyetNjMoiW2JEV6Tc/Ms8XW76I9Dd8w
8NbBrXKWCwAW9i4/VisB34Rr+fNe6LwZ/p5EZpyEgdRhJPEaClX6A26UKNlAOljN
NFpwONbMoNtqwcy2c+c4iGmPoLZOzd7CbV8g1SYfLuKHHbSJXinFpct/+8Z4NZNR
asNlBBUsnI0Ou/o68F5wknU+zpWyKiAKMbqyDhwsqoV0ZAgZ9bDaQzEo6OGZIwQu
J+Inlnn/ZYZFSTkkhg2xth6WfTsc2O95WESnZ+4AcGKaddF/tGQGRdKwFUoLtIDX
SL4+R+xVmFlPJiDXOxhUchBeA33ovsv/9BQNTYH+hl2JPCChjeieZ7lkcJ61snvh
nZtfANtRIoi3MrUUhte2QpD63ur61n8Tf8Nrt6dK9ayq3bym0Zn4jnLPnAtTiUOb
MQpUywYuNq4SGB1GDWp2ZCjKfF309qSHnSk+8jj+EVMUCeTiLeHT+EmhA43vBmn3
gNE+Jwl4/nv3wY/1VNWZ4zbIFiqaHi5mRdIU8pRU5l9ljXm7Vn9D0E1Qel8Ig5gV
wW8WStddhoWqvZJrybIJPge+ondBdLXVsjBsm5fIjbkQCf8pdzdS07BC+HhC0PcL
8Le6daQALesjXGa19DeSla5tDrRDMZIrq0flWYWuGHn/xwLsU2yE8tVCgst9gPOA
OUT0F0QZ747fNSyFs5+N/iA3LqHfa5V88mQUOYPBym/hL2HAGYABlhg31WrCEtMP
9LXdGWr1q1tupnshyNAtiBJKhYRCFi62C8g5JkoCm/Kvrzt6JrnH+LERPawJaq23
8KFyfaIQ1t9zzKQJYHV9uiR2bcpwucAZ2uau/FwHYTe50k/ZrBDrNi41edXo6mBC
8Ok661i19Bx5NNzXb/vsq+HULW+hClREH4H/W1Sk6wy2LduS9VzE0nfcGf/Gf5Ko
h0/gmY31tO38FwOi5609p/xXDNLg16yjzX7zOwVWMaft4kiKlrnOmUwtaus2reYw
1/g1kAvfdHpqv5A3HqkYVIrsJNwojx4+YWttMF8IAJLLOifcGY1o2uvjhPHeQ/uW
JbSQVe4qem+T3DkJy46r6AHOPQnFivkIaMGhY3l1g5Im5G8Ck/0uRWjniSKsWKgA
wA0M8bZQgbzCkJZSllhvS+KOlUP91W3YbyuapCwmjNZkZ/Rp8ucha0Hm1IU8bfrm
A+23T4b+89e0D1cNhT+N77oZAIjWqvvbwpPW2qH1xgals0A4FQGIWRL8rA1Pvn3A
BL0dt5QMEMJWgZ1jrDrUJrLmmKA9fEKE+n/paiMnmeBe75PYs4UxfPbtJLLc6C/x
qR8aVGd5L1QHPF5H8ZOdQTHGHTkaCQRIEfcgxOFNruJJzyNH3Q0IcyszSFD3xh5M
KrJQBxMlA9/QnBMgdNsYXl1YCJxCpgACyVfMyBJFUYMg9JifelaBe5pC1uSvoILr
etoGYweur/27Wb8M/H46/aYk98sHqwZ9+9N5J2tbJ/z46yXXGDAgFGxuNMOBpi4O
0v36rr0w3Ks68srez0+OLhFEm+43Mdam8BaahC1U6ENIpUMnBrMrYDnzGnXqbUsa
HeqG3Zk2OvyGfbca+Mqr9W5ariJRybIoIhhMuTB9EvEXTMdeJuHH03hkvGKad15m
UbpjxAvCiBHutl2R9PuSU3nqgFZzuB24jXJXXvSNAk9GAkhMCBLPD7T9xxRx/LoX
6wSfQTwAHfPI5dCvZgpQz6G0CeInYMgownScO/hM5jXjhihXtAThI+sef6vWVkjl
YC9RKXyX77QmSwTCxAxxYlFrg7AtDhjRikLh7Mhd7B8oJuNZujkEA3vK1TmXtpK/
aJIPMF5GTJzk9mG9Zj6GlJ649lZFH34NS0j5zfgKHNkm9p4x4gpMRojfN+SmSl5A
VBy9I5whJfRtFje2U+z2Ucwzy1EFp4gcP5xY3zp7hh2M4QXYw+n0gYsbx8PVCT/g
AMqa8v3Se4qtVA/oqZRYs6T1E3e5IxR1WkDtGdVhktCJLoHFoBtBp/mkpdpgJfto
iMfaxhozAhINOfInCtwEqS5koXL6wlyy27zuvQRN21PRHQu+w5Qs2ybFxhgbrY/b
GAkaVlA/bkMHTJDPl4yjugnFRTFn4c/OkDntWDiR5VpnPWRd7rPA2YT7QeoKga2E
4dOv8/OTwVHIRF9VAF/IQNELqDBaIajbOT9fbhD/R6cjAzYHxpiazSjmx+eu48mD
ass/SkCi+WNsJnEN6cmHh9JCRGe7zfnaZG1M6DU/BG+jnMGlUZ1MtpVMVz2Ea63S
5ynoaWfzgf2bDlD9NeARp2IEtz90/1uamhKkDijT6bHoIgmjbGM+aFT7xh7qdGkk
a/RvjzKz0l5cvskrYZ60O1Rmq9Qe0x9mEB+8ixvWnLZ+1PGIskSWOdhwREGV5MPC
IP7lnjaoyjmciFG4ufWabODtq8rpdo347evDWMCkexFfXXa6omkxB0Fs2HinHFcO
r0ZsGnSVFOIf6PBwNd0TKghZAEiJHbBTotMw0841eSUyKPGr/BhMM4pkIlWUlR9A
1qxPlheRVsNSB9eF049IxiHBlLJAirAtZ4QXvxxFYVtoTpIInzi/nIl07Wvae6Zs
5s/AfuvQOaxYhdeGH+CO7Ol6SxA6EVJDqNszatmI5x+7H3U1l3cMcUR6njcUixzY
IAZeCRAuL3TgvxRm3GYlcbjhWvUbzwE1vzTYhcwdcBKsvsNdez5bM7bAm5O/Ie6w
f+DyFp1LW/He/1gUicVDRSuQHjOQUZER7lzfdOlAEfEJteT+Sz5Lyj6uxsDwa2LD
1QrJ4NX7opaRKWzqt0WM5o6KMdwgv+LkjxlwBIcoaxd1P4bBLLnXFICp+CcgfQQ9
t7JHm2yq3ZkHDPdv9CxoPTsC27vPNz/LbesyOtM1tbK0a8ENqUO1cko4LoPamfnX
5OsSjXkDhKm3UcNwrDEVXU4bKgsDiaTZjDc5oEhKL4auskD2w8gq6akcHRM/m6GY
AGw73BD9JjwBiIhU/UNfP1BBIsxabtEMfmBpCAbvHf34xj609fkY4XcNJK1IIUhe
Dnzhg7zmp2UBoP/bnNtRO0iKS0Bq3FugLz2JfWjjyVaiPoAJwDYCG9SJSuAJBN6S
IMKt4/p+9nRwHdQMKdUb83sU63ajEYo2gwFwd3BjJx/3Cxf7W6fAMeGcuiA5EqMI
596b6tR/EHGtBHe+aniESoLQzc0kcZU+bS3Xh944uwukq+al0MPIOrxyze0CBx+Z
BscDhkhGYoHnRfngexgKydBM9suAJEt/Pt1fKdYgZJwR3NVjeJj+JZh00BRCs5oi
Z9U5EHXrSlbLwzOBakS/qby3AjY0YvggqgyjTzgUhTMaYH4odSAbdCCaKajShEme
564gizRcIkE+Dv22lRAUORdZIkio4pYL4rSd/CHcK7LmFF2culxx/pd5CKrjTswB
Qx8daoVCaeyHEXg8y99hXGX+xSxZ2jPghM6wNVYNxwJEiG5mkPMBDA+wz6vVxZAX
pQ5qrL0Uf2ZDLqGHntlhqWOwO6ssPD1bA4RBqj1zraVnAV3mani7Oj/Z9APEkQlc
h0LwqOfNJN7u8lbYZ3rEvFTBzFKdVir1DCl7vI0I7LMP8Oay0FWRIdCNUvpFujN8
/PmCeIRvfvHogu/Q1OroqzO/iIkj8R3aOYUkbjdsDHZy7tmQrtzVmoK+cv0sCpJk
oB+5SG/yvCc6ZE+HByq+N6Eq7KWwNBlQPV8Uos4ymea4WV1ngIJKCqgYMzRQssgw
KA92/m8+3ujDwCZu7HC88pNuLzMEPIQJUs89zs4M351kdJ5dqELI9jdj+Q2btcgl
43wLQ2g1u75CxPiq0XlWqykMSDAS01Lz1+msyOYYm/gjsVjBfmCCSTr8D75Rc+SB
GCtLpeGzWyj0NtAPZTD782viT4sZeVVJkktOiTfweVV84ovhxfGNXRgaghqD5cyS
oSgycCBoxZMrH/Z1Xyry6s1X7y55f0WioBCIOQiz4j1l13Ml88bptSL1oQUUzUtx
QSi/eALRekMcDcjbdouGyPNi9qMr1L0UcevQxQGpenj8pG9CPP4mKpgwfUlf3MTs
doFvnT+rZffu5+j1v21prmviRHJ0GH+MLJS+cKueWWfHOv27XmFEepSXhjSYLb/Q
z5dh0waGhD8IxNXSGXHLQjd2GcVEgyNN4YBpnh3iaMEmuStJTIdqdXdAK1rbYcpk
MwHiy0gThVGYQdk1G0+NtOPjsImtxgseoyl44T1yoGPgJjgxNTgBHHxhd77B83NS
TTy9pJC//cWno2gRVdE5nCGjL8b/qmG58icComyxKD3ja5sT0EwJYMlqslupc3eJ
BaCiruvo4lJH/dJTD/RDYYIKH720tjI4RZ0FSYnwwQlHUr+Y22Z5jyE00oClyBhO
R5OzZc/1etBzhHiju5g44hJiF0esd9+P8Tcx/DbtQViT/A+7eVgyJ6YZDGFJK6BZ
asFfsa2X64zVlasQANnR2zdGZa6gFf9/S/52fB4Dqhglm2uNBdJ8hEbL3Z0BtSqK
MQ48VMN/M87GZfTc31em4p4Rc/uMKnqWp9JE3EsnujZNKKtDRB6Ml4liIBJoHbBh
CqdRFl6q/kfOjh3fnEjfsuivNNHU4Lq6eWmHWf2i+i3Lr9TKGokWUrLBZLzQlISq
DB0uersDiSQFY5uzMmTgjiImhn7FtJlJMeTH9cxUCODQU+fiJZqGMNsTpRIdNf7G
OgVSH0LkDzaBeeNemBWzR+2D8hDGEVqVHOuSNXYz+jBeeqzZ/WXtDvHkSWU03p85
iw1miLQjjRP1bE6a7nGbQpsYlAKokYVaakCKGIXq3QreUIOfbxy4BlyJUahBpte5
EpGYJzIMCJ+zm+IXkTyxNLdCEjq+VCQ8wg8oh/o5ApLFt2Es7dCCVdIqw9QoSOXP
fz+pQFEJhlPprawZ1D365M44SnslFHU5LjrbMob0hBt7Hq3IUzg3/1FdL0ghiBqU
NI1cxQw+TGj02LNwEUpJa1py5tXBgM5z1WJQJb2PIizK+4x6scYkqQvLbqsC2Gow
MhuAlSHIy1l7apUYL+LOcfpfjcqo9LTpfM+D62s2BCuulBo7DYnK3PrA7jjAD/qM
KNdJjkMGrIThdfruUT9XnFqtDGPKV5vM3kodeAFD8mITyY8B1G6zgW2yIkLCK6zC
ZGwqT+oTxbq7eSlCvrOjwwVC+V6ZyO2rupR8Hy2CASDt+4kdpTPReYuWa6fs14NE
4AmQTIbVjfAx11Scs42vYZHcaEZHTYnzUGmYN6zauTJVKT+wZkfHomdxAszDkoXt
mprvlze+YyGp8SZZZE1RH4coiwK4HLRU3ZRqdMqKRmsCCk91wd1AuspJcoO2t6uh
v5b6rq66bc5qmWyRbacOKMVNXf7O58EH7n5kbxRlGZo0eEpcwqZZQR40gr/Xw57E
xsgo0vcEdaXf2w61ldHd57War8CfQ04EaNpeUOxBh/+2UVrN+elQhWmlbMPTYDdo
q33n5+ZEXd0qOz5mh59xdWvnBCTg0Bh8lILw8sZEnwIrvb36BRAa5hOHmyD4u/i+
p46t/yAz29Qsk326LEWYUVto+nhChUXhvmrXwCudgl/DA+RNv+CrBdrdFA1Eu8jB
QeODdMZq4dcVBf1RMQmnGLSwqLHnY8ReYEskncBsp0Ql+aQQ3wPlVFVVcUnwOZ4v
kGMnEWe9EYlyBWfC6PIBUtc3g61Lg2QTCFpkWXWTsgZYXy+8MEmeKgR/ORVIEjCx
xfJc7ker7HyLP8FRPTsuxHBggykUe1gWrIFhck7G/mZNLjHJfSXAySoaYpOImnC3
syW/ZFWFZuiug+6KjAdUugtapVym5O9yAmM0WFtlr1NA2JU59r8OBh+f7XX0TwG6
jC+zZxE0cR1bEygNlw4UfWGSSuz4juUmzorNKV4x4mF2QhHvA6jeOXnVseVIr3HQ
fX8b6PAyVoKv9yGJTHudpMfOqxHQRn+8xfx4KZqIKWArhbZpEY/o2XETKEP5MnaG
mqJoJWFyZZGLFjY3B3StKqBZkiVcsWBJ5wDioMX/0hrNjfe6M5RiPxdtE0PXftLi
Rom50SuNlnVWjWIuNqYhqilNAErxYD3fJSzflpKY39MfuMvJw8t31YKFssWIuCS6
avktbe7U5zWJJmxAyBWhAkwvV40AvtfMSuuvrLDWpjeYiKVEZpgDfAsK9xOrjn3g
OVRpomsR4IZ/k8OELS5UtoSD0idujuyVvcAQDcC2mCsIi/VqPJdm+H7Bv1WhBk7z
j7GPVKhIzNET61TnDTJe4I2gOKyn2HSSKr0m93mrqwwpGDb2UZlfboz2Tw7e51a/
xLJEzSl1BukWd3GSks8ffKgrKDcKd8QuDpKpCRCzRW9Sq8gQpQU0tRlAeVYdaSqr
QvLqwrbI6JVR1yyIUxOvWT8htOjpNgOZePJ+855Nu1yhxfLO1A9AZoMzgbwwS4HU
0BiUeDYI42j2XUOrABqNP9iy98S6dXlsrXF1Xv1NHSfUqWJlAlcF795+peB7sf71
7u4TfVw08gaJ633d2polDLpw9i668tEgmI56N9ZqchTGLxzCdruMZAnf3gB/utbj
A6nhmvFOMA8Da5+jBeINBXvEJm6mbepXbFvaSpuaDw2Ao8cRorsh48QCRFeA4ORK
JrvzsGwkEI8fLCW0LF+zpOkP/MJaqNH6VFehpmRkHdjBVEUOMs6v1yMT5ZFl0L7V
AfJOgfbpI8v/bK24agyzevOvL34oiqfhkY2JSvtvnPkm4CEzuryfK4udi7/s5bH5
rjV3ZORaQaD93Ql7dKMuI77ylXjbvULTzI8HRaYumptw4nYqWITFPTD7OJcIbLuD
gX/i6QRmjHkiBzfibnQUdC4mMYZe9WfNZ52WdJWcG2hfL9liXakgbNXX56vD/Od/
Bp2sft15Lf1gnu3K9aATxQ1bsNzdcgLVCWCF6o4L2lBV4dTBB6yqnTGQpg5DlJLO
YqG6csLjSgrUixbdnbeUOo1QPPT+ZLunvCPzh6awJ20W193j5Jgb6+bFbBnoZq3+
OD5zDpOHgKyhlApsu9qZoGR0VAjNZcNfH+d1URwK100GY9nBFysJfk60i/SH/Pnm
Or0I9uchgfBgXAvtSjpBtSeuAq4YgIxmNbIuus/8ZSGoPvOVJDCfuIrIdqE60d0w
Le40KXA7Wq3LwvtAsckAiADZB5aOV4NXikHJs++7krB5u+DpcZtJaHdUb4qKyhAp
kODkd4fpSO0Q8/Eei2WYkqIYtOAMzC8/pUFmSkRz0mcYZtDqkRI3u1Hjb/bsZMUS
itRlalE8VrbB6baxrrqB2zqbKfq9OoB1vMdm1uUMJ5fcvpo2pk1owdyjA2yglLGm
p0FT1JOkvtwL8MXGCQCMvDjZ+fjs9xuBXTMwYT1ghlqN1Uf25ATluiXiINj+CT0L
/F8V0xBwLkQ7SvS+ue5uWOAqgiLcskOQXdAAa34armVHY/qzmNcbRoS7XdbNbNRB
rtjI846zcMyn9GlWPheFV/dak/mQ/NuFhrNkR05DCW8Q9YPbKJ7jxh2ULGE7H/nq
EprQYIzy6ehuswMSDho6xHWv+ZRFy+HU2mX8p5L+8MZh7nyNLymDmfdH4GlFdbci
9s/l8quz+VAXAVwesu0/DsvJ5Hk2EsttNmj5U72unCMtBM7YFYupsaaBertRCNT3
6qcj475Jo7t3+NMB0uwBNadCH/aWhHrE73/2PnzMX9CYG/88AtFm5WVKC0u/a4Nn
o6ubVToQMv554qqPBG1P5rVtK+JHBluLgW46C8inSeY3MCunfvpDlQopT+E49moQ
vQAo+2BVIKhmefO9I4+TEAi1llel8MA+2IXRSVs+MYCcPaTawwaN0KEEQ8D1cRE6
iKSznJv2pfgOibzJjpsPLEud3zOGYcR/MyLpgsql1f2ZpbHBxWfChvIbVNYlQr+l
pk+EjxpTI4YBIXQ3PqboZiaxD813okt0P0nnuM2HVOySdtTygPX+8zHo/g+EoHln
Q8wfq32bG/vNWcROQIQ9QDVcjpADBZsJU0g3Yk+viNZvf0CRieJNs9mxcDQTXaUr
lBM3hJ9a93Z1hAYF9higM8fmFgS37+u9voWBqK1tzmnU/WIVFnV0Gn7WSpji0ZNh
ZNML1E/4bVqjZdpmsVI40NrmOMH2s5R7AQtxoHO0ZD/JSr6BD6kOo1zwX5UIqeyH
wfJ4CyRCdawMwelsx1WpBwEcvSxvQA+H6Co/7WGDNyhiDrcYnzttAMbP+ym51WHh
r+Qznr0nkVdxLR5vVzYWNtxm/m30Jv40XPTlHvoyaghOxuxZZsrViL2G6w/fM1eJ
DnJUyPM+pF1vJAb9A4xUBaRNa3uoTlKOKbtkbPuMmphimvw8P1tBojA1OZFx36Nf
h0VwH7zu0Ze1uAkPuz59m+N+k49ViEnuKrmf8aM/cbdPDwM0b97KfP9LkpLKn/Il
P2eRx8g8Q38OtoNI7ekOFPfB3KD2mbszM3wtZlZ9VwxcBcQA7A2jC/6fU6VBIax4
VUHSFTvMH4PV2omgRywDffPRu4YwRqDM5xvKcw2KliMsdTTtUv6LCMiwbDMDuHi6
RAgkW2ieR/HvbB2+s+194xqVvwsmvLOOteaZyeJt0dTQ8xSf82of0TpVu/+gmpfj
OPSdj5GUcRyFPb1XZH0DuPlBAFOSI25Ja/lri5Xui51nuRyyzGjigUuB2+hSwqWD
Aj6ZnN2/8P8J9/QWPgIagF/5egz/7gQ5Zzq1hmKFPnLhGAqvKnUo6cPHHdaGsSZa
cI5ZIXu6FCWbN7dQXA7wNna2cYi+0AIaQ0UnwzQ8e9HuhpH47wts44KfWpiynYbz
WiwI3lrDAicD5LgEv6gnoho133ztKNq8Rnim8Dd6WdhaEbJ0w//fAJz/1Qbie/Ka
Ntg67o/O1uF8QLPraW0225BE0BuUMZDmOA2o0nkTooHgluhxviiQERIqown6aHDh
4nmEoZSeFjLmRkdy1TAgNXqgkG9F2uOfHVzMKn0DeqF8Ge8z2ILNP1Hdh9ZRccHa
BOCCMnFXjZSbqDgyWJweQdsEWPzV9iJAWz7m4fVvtYAFAfeE13blVUwxd0XrjRh7
AAgfNolqwpgpjRmQY5/4M75ycdYBX2LI1RMZRtXvQlnqcZZN+W0WHXGllK5Izr9x
D8rgIYEtoBnY7EdAkrUipZ4UHbDuceTMNTbQRJ1E+zvP47OcbqH6+abmijwLQg/z
i4TdaVs7GOcesb9JqPFbX0icz1g7yaPmD4G5ZtGymjxx3PYKCvC+douE3oI2idVa
CvaMkQzIbPqhEzoyIjp/0Uvxd0dCwVeDrrnhXh5A2qRJx+IcVGx4MHheaLVWxIzS
q+vCYpG4mS6F351jO/4Q7iSuxSz+cxzMK6hdoFTK37q5qUkgWXDAf3OXKQE/s3IX
tk2JXYTzSSEXlPtgq6ln0btTlifd7v1QtVSPKHUtQFDk7HZgI/2tYbNagiptmbbh
oGT2zdAf90OsqdHwpvkYONFB7cqNNOF+Qo7/4eOdDg7cQhta8Adks3GK2BX5uUtI
gtz8kIHw5/wPaxmrZEosFWOnncXy4BVFvz0QutSlkyCB8LW4DLqRcfFamZphQisu
Xfagvn1DYkF4isjHS0cCNs2V3t5sWLG5T4e+XDy8K71qIDiYZ3vN7ECFxzu2Yrqc
+np4d24e7/gplQYOkFg8B/KfE7daMYZLcWGxbTng3BpK9CqTRV2yr0y3zF+MjoX9
iJ7e4OMtSCsXykpzET+mVUZ7VvjDvQ+LNCAG7Jz8bkYFIIxMKJ1ti0lDJBC+XXCj
usM0ypLLaBP+5k7HZE2hNY0nQn8sZaqjcp++bL5WIFIt7IDaOW+7h9LNIjhyGY1D
FbA8RoSPZl6li9RAV5MeDAJqvZEK76fmElEQx1U4ygZhyOS7YcLteEgT5+JVXmf5
YpZdUEvpnmUikBZOMvGH6ueHjVoC51Mjk+zPw1Qe1KQc06e/I9AZMi6LHOqUbpLU
UMOirIZbnE9hIg21rZA1+vELId7eCp0IHqwY479hfKMTgc3LIW5DVchRqTbyqpGe
frCnZn/QpzXulr0i1zQzicxq+nN7RKyCMUrRl6IsciG18BJRFHXF7grYHZMA1J9v
+IRD27oSvY9Jg+O0slRJvJgtvOWGOZz8+454kAj44S7YLrALbacxVCGZqmK73Me4
/RlfmzhI0Lkt8/yuFT+gJehNTxoMURmVwohB4rO6fekI+19MHnxX4I0sG2lqWuBK
ZTfEDAtXKXTcFKqi5xhyY6TqWYbFoej+kqvphF50l+rSzLW/FZb7y+XYGqo9+d7R
3zPfAfpm7omF8gS4STTd6tOfgvs9jc+ckwSumYatd2A6WCRsLm6+wzzrwW2qeqY5
V8hFEaPvNjG3+6Mlk1ErDhXoRChEpu+e7HmplVGrlt3u9Y2P7nLqSuH13hGu/3YY
ElvRThxwpWuTS8QAxP31LuKEEaLhg4tIdlRs7etwLhbV83LKmOt09K/XBF5pIAXK
HWUOdGWazPwWza0g1JxD56fvz4htUpGxMe9b8304XoDzYbUgFjzjNXWG1+v6OvQn
cHkte6OQywe6qIFPM9vlJfL51g3/wgTCHQdXzXQ2kuiqwxcBIK0GO7bERwzPV03C
rK6BQCi/I+JqdlSQ+EqBi5YFGgZNPamA1gAYyG3d62RzwIwi9H3rnMXjXQqNdUQw
Nlw73//0qfuts2aAeosqIeavbPhyKrJ0Lbicbf+vY2+1e0+Zzdn3km0ProfgVXi2
UKIgJ/YisoD/f2IsU+qQ7Yq12+ZzqYV2AdNaznTYyWDMh4ODvRBfh1UDupxTIMje
uCFpe/7LuY2WEAVsChphBYOnkZ1T6rSgux3uAYkT+IKtc1uIMYrS/wFK+bOVvBbs
Xv4zGEnOiCP9wIoIdXDEUlAiTQ1OJVaPiouB1mM2f4WBLwFUE3aNdh7mjayCbkU7
TVdLkQST/J7p/WX33wmOfxKzyjdgpr9idLTl/QHFodYFDl2PYw5W2AgQ30Qw5dJq
no1kfNobZRuxmWErJUzh7o07+IIUaaiJmikRvCqc2pHbwGrU3v+jMSUa8haWg1TN
Vsub+9LjSKVKoaEhgrHnVd5KFPssZwkQteDcVrK5JqGVuvtJZqkwnhW5LfJZTgA7
ZSMphN+ktYV4sr8LBN/qxjVjWPyf3PDC59v7lwaBlJdjXF35IYmrhgPt2Ha0NfSb
HU8JRSmfYOcUPLwNpKIfEVA7Oj3k+oXrMaSFU+s/CtSBf1uHUljsxcaO+hLxdcpl
y1IysgGidmM8nTAOW5oetODMFJZ7JvLWRbdfJgXn6QSyM8RGa3pHucBioXflU259
HmX3io1NrlpFiKfYzfI24/BHzkGoE1uT7jIEB2nGArXz+q2xUvQfJu42B6Vo6kYL
Yu3zxEcXBEh6AQzXhtUJO7yN6TY6mpU4kILjyhnXq/UwKB1WxhKxKY854A8npagY
qo0Env0JtlprKMDK9gk7q3l8VLyMnhL5LcG491HarO9kdc1LGiIrK39lYLAe67yH
XJI4Rzjc0PyF5I5W7aftN/7Ad08VCp4svciFrolZMTsH52yFjQ57+y106QotBIXQ
W44YXLh/w54np3FzCgodw3TXIIHF+IAesDAzKz1ErCqbA9H05fCKUoQJFXiZr/Fu
Vmw7HUCsNT1ilPMtgtXNJmz5rl2fwVZHgKe19wd8PO3heZ9uOZQr1NX/4ZyvrGn5
q0Y4vJOIaSsle28UOZgjGCKnw6hS7iXObFcbbMOKJkgLy/11zLnFl4K/Q+uRgLNV
CoaONTixDKzACLOuNUvIxXZ5roCRynRjgUbgjAitY033txeq6X+WLrwkCjgwjRTX
v9Ni+nu4k2Ct9IapBlFrxNXdtX7K6n8IBsqQjynDiHLBIifBUdJoYPN6IZ8hGYUt
XNF+KeLc2La4aat+nvrLqfSz2dhRhyiRCJfCTnudLASQRikXtPV5sUnpm5cfo+09
+MuhOSt80/R5VppPPMeVcx1WrEdjXuZBFVO68zh5p+zE8FCpmJetiMIB/3WKRebX
FL1EhraiFkMTlFyJYH0FUXAck/GcWHKw5dVUI6hVK0KkPzhr6dlIpnPqh+rm/8AT
FfPX8nsmV8l7E1Oteu9gDaogoXMClaIQggO2FLeo42VtnX5csakve6Wremhf9pB9
jvVaOSTVk/6FhlXLc9g6J5HkJj4piDKYyZNoieP+V3QJJDgxdXZ4wYWaQNEiAFUw
XIa8f3B6c7P9Lyy2F7Mp8fxcJBZLC8kiWvf5XCjrcnyeRX0f7me1AnnQYZ1Z8gCD
lUV16T7b8rNJ2U7hAkViSbkivQUJ1ouqwcLjVp82Bv66hAPHjgavY7KyFrKc9NJ1
klGt2aO+cQVPLgYeLgJPhTmBXEahpHnJV9RsTaKYffjOqEcTCXJ9juNe6xQbyeSp
lQr9798iyajutvIyuo7oMhb+3qRaKgOpQEL+aIzLELXM5c+yNeZCoNuFlXT6mk16
YR38Q27Z146sHYDZ03W5IKMWMZwRuqgYpEImRPXV55npTDxGRDKEhpMKslpR25Mw
OHVHkl8qeiV/InCrqjn81XpOEkGb88gWI1bJZNpUssuj0mnd6/DUQC05VxZwwELV
pD5YUNncDvnZpT1xZjhs86I8B5wluMG1rEveJr6kB4rEndB72HxQGDx01jDwBj9Z
R33/OYSKTx/4j6AJr/8opUetoQ5f3uooGoJqn1J4nvu1VtanaDwGAIYMbGOtw76F
epNvLi84LlmnMUSs+TreU5N6e6A/d1pwsVWFumJhAKTSKDkDFIEPSpucUiQFbZhe
v4QaWXNtQRm5PEIkAbZR7gxVDGlq32SKQ7iiWk3Dh0HffiRdGSHq4LRckcxk5tIc
2m7brSbYhPW0n2nQDCEP2S9f3jXCCa4gbqhFlWl3D6u7/bwkT5C5MbM+o3Vmi28Q
pQIVn+rIVZwvn7a62oUdxrTrNoI4FpU16Up/6LbhnpkSR0Mc8VemT5lEMuEbfhvW
P7RxqtaVU4ZMIIp3/eqm45AmowLOGO//PMc0iabCvSexaQTE+FZlx0EbeDiqbPlI
TIe2hAih+1E87q4/kXGDl0cZDDG8VvnjWsC0t4J0SVZ9d5VBlERXH/qoP6OZqG0n
5wDtwqedVJ7PGCAGfTo2crnuFus7jcFsJCeeEhCbkGjg2Dct3n9MAT3uFK00HNgg
zvjRBkOQQrrCXEzxBCy0QMHW1RI9sk8Z9Y6KYnSnwHe2XkGGm+buMli/G5hqAXva
aiR2iwvmztRzamnuXXL0YJw+KkWRyYj2fafwaOPAx2Smr7FgAHCQDcWl2JJDLP4b
CjEHw2v0EQZ+Bnw9MdzUUO5Iz6GFi+2nbTinGe8aGeBpY2Cyj+bYLHP46BMx6rkC
Wyb5xi9uHclILNoPmmWcGMNYLSNMGIo2m/gIN9TNN0REFMdnRIBTaPp7jjR7e38o
pL2B2xVQ8cRh6wTt6gq3bufL/0kYpb44//s4n4Do4Abv3SXXIR1H0hFw9uzo4pPL
ZnfDAeuo8XO7lXBGNRL2svMSmK1tRykBmshiW2B1nfCkw4Kvy4xrPQs91M9Onnf/
M82EL2EvTL80JHq7CDqnPDrTe0ToAG08yMdbEkSxwamxR+TNmV9rKUKkSv8UwWRX
KibjdVeopVVLtynr+jUP7/u0pW2wEisgjnR5rIOXixAP2JVRjmKnfonuwgY80rF8
XlRIdLODA9k9ezoq2CNqjvvy8qw6VRSbgkNbOzphiLhWzxtk08yn09FocrnFTr6s
MfubZQTulFHe9634e72Mkk9M6K/jqHpQrVmfaa70MTmBe0MUO7mUjqnBRYFlAZ/Z
aU5/QGlQeVyVYIm5G1YTOOGFkAcLhhw2Se/THJIdm4jNNzgY8XzcFRw1yFZ89Fr8
VyhPhnaHuS3MTgbh2G0nfutgvbHveFWHq74D6CjQMNm/LVe95DBQHTb6tQNo8JE0
t32lTInCv68mDkMt8cbBexXDdDviEbRL8tt8fCz5eyYusEedq9GJ6tKPUkx0Tvht
26WsXG73u+lIiicsuafX5jxYTg2A0Assty3eEw8rTFla/BChZ02SNtyGUx6UZD7z
dR9i90q8ZgMYyJMGGMVPauM8e0nv5QcH+5FctOsdSgjdp/GOqGymu4nWrgSZ40rv
167df8o0o3+UGRQ5KvzGQFMkNJQJNq6ocmcTCQ0647CWGFpUySi74fz8fUx5qQ/k
n36ksArv7NgmE0W/sAnbt3355YvTHkUWUSwEWU7gk6y6UsqDeiR76Tba7eq7tr7K
9We+ZB74xnWklgV6P0t7cQgrOjRNem/9MSFxv4FvSIiR4ZStFe1skkfJpXI95bhe
XEXO37RSWzV0FP+JIeSa4ufDdmvS6wJnsyUYwQ83h8GO8qGmjIey2ohx2NQkEFf9
9rJK/3m7ObekwNkC/9P1L6UD/xjokHRzNISuJyqyDkcYQ9n54Yq4QYajarY74zqg
WK2abQ8qqMeu0Sm/HP3Oqh2nYkCHtgqmnXjR9TRUhdGDh2OlUe0L0lHGq8Ln/fCY
q1Ghn+ARnQX/OeZzWm0hktIWHDuWdOLqRslmmDfSlD9o7GBhqcKCjihIdD4mqyzK
w5T8oXiRqeu26OReVi+NbZOf78FhYLhYN53/gQ4gqyYGJI55VqVLeDHi5mJJX6I9
YhdZNCFrvG+ZcKDGJMdaWvgoSBv9dLkU4TORLe9//EZvOBxERObeyWJB3LNUxwp+
stRrXdLXKnzyNnp2uW7cmnBTqEJ9AiTxyoehG/k0XXNyRfTqPI3gmt9ZE4Nm8ug/
qa+bCk67rXXtr2IkDkGMBvLXsOGD2Xt8GK/AivDnQydopFj8XkufeNmKyCRdcPDk
CRbETcEwRzajb9zEO75V4K4rHW2AO/eY4qCPyHY9G1JkfBQw2O6oG7ARURtOO3mB
Eur49gJoRbFbpsPVx/uOuFAyp7BqutX1lfK6+L6ulaRviGbxo8oZD6NPfqE+g6W9
L38DEoOmeMc2hD0J3tI3uDwA/yzvuq+BpEuGkiq2Ii1Ja2HucHpVNaanGhZTD9Df
zRFGuJ4WHxLAtzp+uFXWYD1Xr/K4Bmm+UDiK3cWs3UElQWMPbHvKE5JhDflWz2MK
VvUe0pHDhY5zgUdUUogA7S7Zl+3ru6BZ6ZOSeaom39ZKJUkQL6998j6FUys18uG6
yItfHz9Lz/NvSwix7p6ENfRSV/i7Qkc3qYelr/GDcuYB7Blzx0H7pHQBIPCiX3RU
AQ9FbGBdDXXdYe8JfYNSm2wdXXR0aCjmFXrYmY8izetGzEDctj38tr2VI8y18MOI
APJlRQb8Im5L5jN36Q+imWLJNIVd+GreU90RfRSd/xjMhbE20+vEbGOKN90pJAsm
6uxnls8408RFuEql1XaG55pfEFhIHJjaC7QMGR3YLxb8eTjzKgq0b2z/wrHBuF3q
rRQjXtdekzRaO3b5pLpahQfZOvOeDeFogL0EUdym0lUnJB4uG+d+nneIUhs22hk4
h17CbJGyAXTJ8+OeSkBZi98twOUf9ZkEJTn6DCIN1TpWgP16rHNt4esi98orUOEH
cyX81N8qzpYq7fWgguRhx6+y8oSbuwZB4hRbFl2+4gGAVmw0ZVoO4GfI9ic9Sash
9Z+ireKvQGED63DlqVArdb6/pbcEqKLclu/qmOwlQVmJcj/T9NvfVhk51HvwaNSb
gyKCK1RPqftMUL+Tm8XgwuZxri8mGz3qFA3Aeiork1spzQcNqOeyMJ95T/sVQAVK
OuKZCJ9Hrklqkt1fKM00dGrKuPGHhOfPvTeJuEw7ItnBEO7wydKJA91BUTDzdMPP
SeL5UU8N6ns211tAFAd96K13GSPE12cEqHJTcSVAAhiocZJfRbPxDg/TZ0l3favf
lmHZIC4SaQI+nRPRT7lgbzE8aO7AUckhiOdJiyGEP0Di+FTQ6sSJK2RaGAyDh77N
+C9ZzvfDbvpaGNtjMjrKIcH3AtbJUL0He81Nk4xPDL8jaLyYqWcitYyOiBs0UOwW
qjujtN1aLXM7txHm93AEorT6Syje+8xEIsRCRMsKOmklBPkJIqTe2U4nXg2mtDYP
+ZqskX6HksZLpimUzq17LyYaxSZNKLtNqM0jCHWyGj2PVRdEG9mLXQVJd1/VNuBH
ZRI5Ur+uDzr2d8OItU3oyu/cdH12iP2lR6AK1/ewbDnCQ9rvDQll0idZ6cjfL0Ah
xmkqKKTe6tj7RV5ipnb6CDRlTFpUvsZUAQuHwe930TcCzjRhpmQGtL0A/WeJ5ZAS
ydl1UbIGw+sv7guBrJMO5C8G2XQA28eUrXXBPg4qZWQaV4OoekdnPSjOalhhrtaF
vuUsghBc+WaKtlWOCOq9C20iuiC6XdWpysghztlG+sh9aXL78uxu+5Tq+yKV8Btc
gu3a0ddQRvQbWtji8uwNhzClXMXiV/VbOG757+7MAiKGqKmKXOSQ+RLDTG5GF6F4
aJxjwRwtjBdZXjkgcbtLfXRYBJyhAuINNXPyWpyppBde4zxKXsDFhb/UPnBHktms
qxQLl6jf1UI/O5S6r7UgVbr+aH270/uoJoFxFdzpuOqkJFtf8siIVKvRu005eSkC
N8axIJcqpm+j2d98aqm0+8cXL06BaY5xkL5EbngwaGJm1g1x3m46KyrgXcIZutTf
G1FoyUHyuRq+iLLMcrDvLMPjWbjelFEDrWwLoXs0xkCJeHCbmurBmLXfpajWTNC7
M/WMU10j8GUyRlrlKv6sMSLD8iggFeeWrm91kmpng0sbqa2qIWqAbPs+QElZlTFj
1eWMFwPJhC4l9ksqjbQ8sAti9lQQilupGlg9DKLgCnWL7OGz4OmCUhO/aBIcvmld
VyiCdj5ENfop65SG3sbSXhb7R4Vi59LdQQqwcV76YmxznDEv9boE9k8euTl9hs2J
jN0GJkR/maDz8h02m1Mx8ADzOQK3Im3wBej5ExHC+SZmYmE+UG1fEAQOq/EiwYd5
8at7/dQFhCpcXKu1Y4c2bvJmRPVBvzX+Y/0WSQ7LJxWACvT1A5k+/wuJvBcQ0kyR
oSiQCKUjSRfDo+dUQKBmJarxSjRXX4HnPHrasr302jHhxbRb548nr1g18a2C0eCM
xbDDmJAnF73mTBqPZWHKqbwS2gdNiuUB/DlBR3Vz58n0I/W/xdeL3kIwFYuoOAV7
WqEtgJ+rjIIEHi2nLOKksCPcminApmMOcmHqEuekusonF9vsmRhgvDFgvzPkjBxl
vBm1sisnarDmv3Qfq3Fl/cbno887Hse8hnsZl6998aCJeUVuYJZYDL97+BLHvyyW
/NWhoDs/HCYtq0YMNM5MLEfT0k5qt+42TnP4/XdwxQelKDgqGCvPCjucy+5WUu9t
10BQ82e8jQby1mWcNkFKCol+Rx/clgUBRMMwQuMbRjA9MYtsDMiiFF3CyNlB0Ign
F5CBaLm5seVsPXRt/QMB3D+SlN17cjrOcGAAjy3vrstUyXN5poTX64b+Q+zGMXDR
NlNwb0KpiG50iNHPxhOxGehRKjXCilX2I9FBIv7XPR5GrryWTOAuRtW3oAaU8QNc
yE+aISym0O5GOFMWJIB2UDNISEUhIxy4l+PiFPVdL0dCNuY8mTWKdNw2olXd+E0c
BQHdtbyrd1rS2gUJerfe3LzzzXlVS4YgZG5yWvTOSYnIyml5iVFqX9u+duXAkE6r
l3kb3OFUNBIEjKRPtbzAJRXMOANZDKvRGWypCvoXSvjt0FBkSudIWqxdb05/Gser
0OQuBw3UT8eYGdPUPqkJhu7gHXozuoqcA/R5fD0tAIlbaQna5pmJczVHpPAP3HNw
/eANly7sxvrwIeZRwpEu6gs9TrIaSUqQqPZTe8BCMdb5YqyeR8cTvTEEBV388N+z
YvyHXIsGLw5j7pa/eBYf2ZC1+2ACmiknGDcRfOdgwQBzWvWjHZxCf8F969YgnaPy
Ej0HwzOvmPuKno0yo3Qza4NeMp/TJeUZn6/IQcW+8BhjOSixn+Ix89Q9FaXbI6gr
JKCRSD5bC9RFi0j/RM20E+cfiH37yFR+KoTsIW2Gbe343y5yOrdizHXrTvnoSM32
mqBHenfx9YrYYwwKz9iAVSKzYTqSCVU9VuCJSYXJkmYvwrxHtW2MfvI0bXNh7JYx
ynpL9yUzW6+VdLOf7r2774fXDaUOApRU4EOcE+F/xDIFG4vPsJgG4ZnP+wghVzYI
++Ere3rZpJ0zxz7pfC7CUDfRGxPXsp5h1aufQYo1sD6i+hkVI6rKfc2N0Q8M50DR
J3PYDgXbhAGbqTOzuNQLw7i5nKP7ueeag7s+BlnyMqynJpuIqK2RcLxbpDK871eG
UUYYC9AtqHU5TjB3Vx2VzSXg4dCnmNmRs/q3tFprNrNovEaKBbwxXdYfWe9MURQB
JrGgOVIb83c6iI4I+vkmZ+LYPBgevC0PyY/VhUg/rOIJDyEMEAX8JPKXpwHV6PZb
9Q3cQ++Du/A21HY68QOZib7iDp1NMQbf4XJArwcjU3qSh21vq543mvZLxXJnLXJ0
kA72FjkbzLavr9+9R83dL16YaGuxiyUKbyVLmU2telCaoWF7sjeHiPG9+DAAj21j
QBK2G8SZjPVt7HFosoFDt/TkstHrHDNgByZYPCEkVVJ2gKg5frO+sPDNAt5JETgn
UdoDWNUKcM0RA85Xk4Nq1HHI/eFYFbnIM8hPQJ7UBQcZZzOG6faaN34Sbi/rEW47
aCzqJ1B4yXJyumpJdVqKXp2fsbzOxRCPeMGLsGJDllPLMGw8+hNCZtRalEUyZajU
sxYROTCwNaKRfe9yWGOAWs50PYZhTwjmHkdXtJCBK0Ta0wRqjAVdfKUFwSLXPJek
pxs9l8zKUcue8ZHDtf5cXlS8+ySQan8PiS2L/hjnYExmmtajHxHoiIgOz211gGKD
ALGLdTCWch83ICLZCWQGxR/XSq3VL5Y81iumkh7VA+xs6FgvaOtrZU0EytWak/+e
CNxwDZQ9vEgogYOfcK5ZOe9y4IwcRRXUHyFtUqEqocRZu+ROq0ylTMlT/uCFvk9p
CzG2wTt8uisuziBeFh0PqQybuy/Dk5refl3PSP5X96yTmOQ22EVzHAHg6MznuMlY
+LfOegkvfhDvTN3Tl076lZR5kbU+RCP+AG8D5NVg6Kjjb20hlvi97UAoZrRUbeju
Xj704PJr4ozUTJixaNNucFL5AwDPyxgvKRNrPJFbFoHGcwspk8lLro+510a0mwhu
Iyq0bIiURrV4uV8d6eVx1b5Dy/rG3xGLAp7/vn19ewRxIG+Vi3ycRgo7XKHzyi8o
ZrFhKa1hwANphFIT2OVWj2dhsDiwuWd1l42MJmixYYuduDCjrJ7MRHhKo9EoCnw9
d3XwVwuUjQfj1esfTuRN7nrw8JUIAZtM3DKXPu7cZS6srQ+vubt8DP75a4ge9Ktr
RaGHJrGxOKcHTa+KfiIuasXjEk6CEfNjNVE79rHQikw2P10QNNv1KoA/QKyowg7c
oIcLmJKlSzGrqDbDeEGqBfsPrBfCRqKtBTnMmN9pzdIqt5bIF7I3vmQMP82JVjoX
L6xro6VXPotLXPcas4514ocATQI95OLMWHKfHiM9bYPsU82bSMg3j0K9mLWW4+tg
Q7Vknq+IYLJYYautfZTg1O31OZtYL4Y9Plp3ozbJhp0MeGB/Qidig7MdqCh2NIeE
JwpeUeyn4uJFa3Y20aHfyMHsJZ1lsWIDtwOtvVSFoTjBq/rHCi+s7cwZrhAyyXkw
uHeOlagWr/NCQ4PgYy2sGGNzHbDVZhJQMfsLdL+ytILEvY+t07CQoNUFnUGyxuDv
jGclTKl36JI+8j2eUW1ELl8Aid22f0UJqbe5yedhvQ2SrnyT688cNYMyxIvU6Jv0
maARMa/goHYY3R5T2OumrBBD01QVIeLIBrMwWJhn47FUGpBYsgV96sD7J4D26up4
oZ8GPAiOutCHZ0K2p3suIBE/KFai6xbF37u3vYDtQrlHZy7KfRKlk+FqIIH11AWQ
r9wnMhZrLhh/Gwyxi1X73+RY5NRNKNHlqM1J4v957Fod5l8CHPDvKL+y7zKsEsgn
xaFvEJZagZ7eTRILfgKM4DSwX6g/PsyodY6oaNRP1DmXNEDRcf5M1QvxWV39/msg
fqwhLd4we2nnq4THfR3NM7QmjXvRa8BIgM53NAFygsMNMdEdnCkRAMeqCEQxXnHw
cHKkPvikJgnmrakg+gQEPClV+TJKianOuRpokb1CorQsGs3WW60Ek2KvDdevBYz9
gcMORXo22V2zCeSx40M4sIKmzmnpMC+RQLbIRmCIwSL5w9Z0iILMGHc6viBmB4Sh
67B1inVDbCZro3AIvf4WIlAVp5sMjk5MfcW5X5HyY9IKboqorlM21pl8/BMq1+ZU
fJRJaTJZxCM8hFjua8965s2LFJvk5Q9xKeImwF3nsvW7PcWGTt/kxB88AwLtM9+a
IdsQlam/XgUn7eSVS1pk+yl+Gha4N2Xy22kVivGuLV7+N6NxFuv1W9gl5ZLsZXsA
vNKb7/V30RWIS5OAn8nVyjxZ+PUhTcr734fb0cJdhu9wmDXhZbE7YS0zLPlt4e56
IXI2wvbUoGwNejnZwqPCaTgJV1IO7/WYH1Ej6qRwfaoosGKcmDY6hzK8IeCBd9Ag
cgIwyzbVXjE7ogz+9mUXxl+NftLEyEkcGKmeNq3QTFVGqlMDbE+WeynvWT/KJMPl
TfqXKdhwCN+29OTaND1OjJTdAuWkByJ4HoF7ud3FQDfu6x2zMBs9ZJ8L/e6aCPr9
3VsHyd4/4yq+Dtp4sT3NKBk3v0fllgR69aDdaplfpPWtSa5xmJEK6f5Q73I6oi7i
yZ8yN51sJtt4upmcQP2XEiGFEyO4ft1C8jR3bTVfMzDZRWbQ15XeQb/QYzOL5KpE
qAuCtOplUF8vUlw/saCGFIoyzvo+pgWcu32G0o1gfJMGjtGZfjw9emrcOv5B/hYA
XnDkFFDEkae2HD8AhHM7U0xsmuAv9knKf3TKWXRNMa2WbZy4l5X/UC5nlSLc8R60
50JTehnHR8akU8wXUl0W8IUyz1HquNqzSNB16X5JHD4dX1zaXXSeGsf7YFP/CGMZ
+coeKc2+8U8cIOSN7Xqtf3ek5mq4IheOwkGNre8ygFKOpGc8BKWSLrl128WcuA5Z
s9mPYO+e2rSQL7MqsruCu0rf/Pt5Tj36QiU3cgCUvMhEd+W2LiQA2eamtTNQk3D/
a2odMZwi5FYHhwT183dhVwjrob/+oTrR/ADxjA1P2mNzdG7q3H6PsRW2I8Icfl3g
jq+mm+fsiBb6E6OFt3PV6kKcGaLakYo+VCFkvmDHw2e4BOnrKhYfnBnMRxWuRP5d
8/qBBU3DK1Z/XE3MvvPgzMl8VTnnBIK1/rS/oc6H75H/F9a3DXb0gXEaHt2f9t9C
/fW1kWBJft/cRIxvT8meZAIKE7YxTxNYdI0ELrOcRxqYgJ7aZB7Hdt59/6Jwv1uM
MAj20RVzKqFG6cZn466jJdqNaORwrBghoBgUwl6ulG1PQ2bNVdViHNStMaUaM74C
1EdqvP8GCH+4Nk7lZKALCFpqPW2ybMFc0q6SbHQ6vFYFanUsKZAB4mQ4OsmOTWbD
+IG9d+XxZDg1EJQ5za0z+MTH+S9gHa+rqLNYTIJ//SSABwEhqxLCxceI+Tipy6C1
TZ7D4Mko4RQbHNoLNa2L9NM8pj+YtsttfkguhFBzqFzkHykNQahg8pUifK1ldYOE
fEmpHBDOfEMuDnBWYlGtONtW1JokAj9nLZ5LLSqVSaVWoBgWzOQ09eX6p/59uv7U
hqg8KUOqng8OK/ogkUwVPzUnEvFnzFDE/IyUXT9JkzgbCawtu+rXS/u4ggUkV4iD
cTUm1q7pXij/Voz8GR3EiOnCZbzjNqT8PbZAM8Dy8eqtb6SSAkuq1THCcFIfVHiP
m6Tf4NvPVbfqkJqv/UY4KdpSuqO7SBt88XJL9PBfy8w3owzoWo3kuRJeVnLi3/Hx
HxFXleNe9hdt8ymVeaJ0dfiG8xAXFtM12Nx8AV1mhw4F9iXgRe5bu31Pelxh/hG9
cT2T4vmCqATaeQuEVM8bieaGQ6Vb2OdwbTRCf3aABHOz9NUjbELxli8nQG/STcmF
nr326660jJtOOwU+4IWai29hm81PBDYw+S9FNac2cStR+9vCG8IPZODH0TR3v92o
I0e8RA1oBw5AA5CRv5aYENoJCnWZ0zas9j83Jxvm+mgyAuTrkFkZYV+0YHGF01C2
Q6gqD16hf9XfCFYAkPBcZCuDBthLktfEYuBQSS2xSl6rbm9/MdBC2AOkarKkqdKj
XXuqPwLWJgkt8OIzDvFV3obBPNcDmNwPPv0BfeCmPVXSCW+7CyY4/2+jtKLfmjQp
rwRGiPiGsIQFGyrmIdmMU5kq/mv1/swsvfxy1eTYsKP/FbZo+MeoQ0wwKuVk+qy4
Kh+WboNjDZXNBTisjkJ+M7wjtgYp9wHqjW0mRKLiO3KGPFlB+m2CxNBWWTGtwt4H
hCNvKrITfkr+W/VYsfwCzEuMktxZEoTlZYn0gYzoZRqcqDK652EsX7P2yJiYDo0C
`protect end_protected