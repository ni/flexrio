`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10080 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/ehEUpUyrMJ5tzBynAl6izHo
hE/NpzDlYOgPzMmQaRb+R5bMclviEqCAQzcvVGHmm9zHg+pHEbH/Jio0DY52LS5H
HHT5cPN89qnaRq4Fuy2jl0U2XWIB90pIhi0X4PRZOIzkyz7/xIgOaltI/2Z7hvYy
NuyljHgYmNvpDo9VS0nTTy2hCnMjHlBrLgolROcxIsv/7Has0uUbL0nAughcNhoW
ZbExoWQildN9BHQEuZ60VkNbjmhT7SNKw5M8UxjpyzTbj8+bzeDAn73HHTJaRwh/
jsTb6o4ONPSSC0vJK5ZMcA5caZBM4P6zqWy0U6LV6NuQAYh1Q9lkm8DRwjh4hk8q
7XGBOuffAjQhLCTb2ORplGH1Wl8+B2QxLuqIanf3D1LC2dkHxdPeFqbC1RfWZkgu
n1Y3FtiML1NLjZ7DBwvtVEWxQBYWPAeoxQIXvMKUg+WK9EIVZvNLq7VyCYQaJueq
gH2tozC/8L+OfhIAC2Dz8r6Bx8FfAsnyWx42w1QjB0lp1dV7hI4SFADHIJ0LBeq/
VFE85P7rm4J0Css0aaysykUQhdEbA4suB/pLGFCdPNrXystt2MWLX4mhACHxQWot
H3MMMR7RSlmgVMYIQnPnEs61MU+G3StAP7ctmRCU+mztQmUMYIGukxoZCgfd+tr+
sAA/zo+ByEquPNNv/+/NRa7C9wsgjb763WZCWEEXajm1BwaCJOOb1SlE0FS4cHC1
IzCzKo3C70oi2kBChGn+gCIE9H/+GxklT85W7Yz+EbM+wdrCoGt6Z7EJgB/IwgDz
cHScFeX8izt05JspCzHGmMmtWiu3dUKRTnU3rvP7bcADVFd2GZQFuZn+yH4zXdR+
xbkIS61ExRGElxi9OmiZq25cQPOpXS2w3J7KegnpQVVBXpuScr1kRweptFrOjNCX
XjBLX0h2E6C6Uz7wzw3YkBsbgfEaBVkdv6c78TCFB6GnRo2+ouwrE/dnofT3G+HX
LVMEZLsNZqO6vAIFimdk5GKmdNRsiHGL94up2Bj0fQMVCPkw+lQeiI0sa2nivIv8
tMitK8udvHVarGywnSa/1BUqk0l7D112+Avi1PPDn2IvV8kBBsrbN6wQLUuiQhzu
/hWra5NvRHJMs3nLCqRjJo2kyqmAqEUdkJ41+i3CZ0zYEcwMt8tKaFTOgXcZnXmI
x9DC8qCJTmOSy5hibmm5QOFqMDXhXIe7qKKsLg+DN2f2kI9fEXg/ubKLTOvFTw+O
UichlMTc0t8N4C85VsuRxkzi8JI8eyaCEh5SMBTnZHmMcxks0u/Ra6Yhwt0qz4d8
PL4w+z9fiBdgnbx1fzMaIciJ/IRRz0LAm+1h3HUQYZHFrigYJ71opXTbz2X4lzl1
4ScP63BCUCXoGNYwrOd75Z3P0rr99qj7t0CcvNQ3AT5VfsAtMQUQ1CaNrEeypWJ1
q5gjKvJ2YgjKARmHpORIJM2F/jlx+sUK3t8QS6J34ODp0RdlFqEEUXcIBJVuw0Z1
SxZSN5iXD3SJS3P88yw8hOSuMDnh81PpXyCMjP/JVNPZkbAFGN8XHZEM6WQnybUw
1tBBDDM0RRMCkR9TOGE5Si6oqqgAvRDBxG9Ksw+bXaCHK5je1vJj1dEg1xx3cjvp
uhoYBnGbnHtYaHvyMH0AGY4jk0udHuQh3X+RYSsEKktzD1gMQTwrEV9Emq4McBUW
qar+o5Ve86okH3sx/9mCBi8akvMClHchTpR8v9rIOJKs4NEpcfe7zo2Kszqx4E3O
EnLMJ8pVEb+AEkaKMHRsmBdN2Z6RJuraURP1RYAyPnSW6dIatCvQEZkk0wmUzpyA
9qhj4JRh5jK/n38bqVLyaaZ6RgQL0IwDkZRurZ4bS8OiBBtlR/vPt8nyRz7XQjOQ
2zwBllpk5xKqqAaJsq7TGE2VDMmtgpWbm3V4C6X874QXATB8pOJnJIrVEVZ/XiTB
6brKysFH6I+lS4f3JXneFF+XL1kOFTOlwl1oXxQI/CXuhAdFhSnp81lGvr23p9O2
YzwUYPvWvN7TiXTIA0JC6M24GTryB1nWq/BRg0fv6njqha8hSShtKpJc5Ymg0Xtk
3Od7f298FgGeBTk1G3Q1/05IggdjEQzjaJZK3UmEciUT6nmMVM4GBFE8mAHcDfcA
fKNufl7Iq20nTsq9RlXvIAE7O0CP89oHqo5/ulEjYFFrFp/39eNZ8MRFqLRu7vrr
f5CPsm7hvDXz55lyeBqNRn/qLhuvTS7z8x1fXbtSaQuZ0lgGk3PLc8uQmNw5Al1U
tKKP9wjAZsjpVktm3X41ON/uoszYrHMmxVoz6VhIXm5iJaoguuVg4PDqR7r0WH0I
IrvjogJmyhxZehHNKlTRWvklbmhGi6Ll7dUv53LkArVcZvQPneSB0OofBQporUiD
0ukaoOy50U4IyvHU23+QHQddE9mnug3xkR5YpGz5UugQ9qDriDcsiyGASyvJM02t
MYo+UNctpxQwMEixXqP/OtJ7s6dEAKqWSLMFyu9gP8HkCofGFOAJWp7AS/0vYzg9
Zb0AIWpf4MnmoffegcigIYRxNxQJFlFABFAzkMbovI1V8/2nDkUNYxAgcF3N8v9y
xkaztzlH9QD56YeWBteW5JW94OnPrFE8CS/Dp3bvzsCZr+k3nVlArnvLbPAeO57l
hzyfoJc3ybl/kGP5dFEoRyCFKH03KZprv1vaM/pO3kpfy7o1Ln/RmQsq2/w9EBB1
iwoTM8L5Itkx8M1Wz1bevMt9mErAZPvjhBC0ce6Uw7rNbFEoRAulgCrV74Nq7fw1
oYm0S0GMCEZSyo4d4TA7NyjqIESWI1GghGktQsHl8OxnZgZg4GlPwa3oFqygu+W5
TBV8wgLKPhcjl+F87MfJuArxnzk7QYQNc7c09ZSNr+jEykeQySXbQrG8dY045tMY
PH5aPZ3gb5mLGbJxxYCSDkAYPqVrGeVQCnlFYqoyA2fOUkFmaA72lvxaXWLt7XQD
mW9GhwxszqcNjhryXTf0YjHhvAFuscv5HNpp/jbvZ2qQob9ioykr60KjiFAaWY0b
CG6GF4S0IGTezxgJnehhan/UCQ+feK5dc3XuOQtL4WN0c+QBlSIXyjPPwOxQohKH
0JH2pKU/4Ks3HFx4Ue5QpYnI2h//+K7pxhk2XuFcXmUzRYtErtGLBBJZyYCLLcpu
l6xsfQz9DDYPt60xnWLyRAy0RNJizbU5njy3nnbURRXyOO1AcwGDCji4QZH9MUz8
8UXhvDYKmo01kFx3IXSksS+Res+ybABARdEf00bEsbO1/GH1b/0NpstAuqdu3Yjs
ZUaABPhN6XOdM5YpVmkk455AlxFGedJ71/IBYH4MYskQzDycTNnSRBlvO9yBpDvR
XfwPVS3rI3/UTQN/JKqUKlHO4Eg0HATiIjHS2uo69lTCJSk1koEzdsM5A2Bgy3RN
KCFb1FG5c2OmsTomTKfaubAsorqGEUNUW+4R0+hdV7Y7MH+0eQi6YmkSVkj5tt39
zvYuC5lQgE2yOh21c+EO9Wyo2aR365Ie0Kx8xGJVJtDlgXFioyuWM+SmWCMvN7go
Iy06UZooTcXe3Rg6/Q9EQERQcCC6yQhIEPtryEerdBWETXsc3GDcCUWrRC2LwDxg
5q9A96zJMGg97QeG4WZlK48+GbfJks5KZxlkOxNPPF1IoIuaOULA/XY7sZs2idf6
bUc0n8DIiKInQGTWpFRYingOB7//psHvhYzqYWcdg6mS63AdYOZExzaV5znhY/59
D47iEknYlDx986ObClr7jL0ijprgKwyFJYtttTlbgaEUTaFjvgnCtfNc1SL1dv7h
vag3GdYF7OuIbyDep2ShxYgEjOqZoHKOJu+avukjzQQfvM0Bw6cbmbTO+rn08reF
ypiH5mWCGhyKK+JI82Xox4shweS7MBWtcEVek6HfWC/yT1Uu4WbRi4HQ7afVdVyQ
Tp0eNLDUlcjUg0UCDU/FMEV3tYRcU4rtk2nQ1dHrBJv+eU5Bg8dnMFIJYxjG6tXH
yMXL8MmpbLaHXUq7FBheR9Tjey64u3dikNv909n2aYJ+GWUYjt2+YRuQ/Cfj3SGy
WafLESYufQdGTPnyRX2DR4TOGUUFeeuUYtGCX1d/GeKQF6pUa3aSzMCVqMmW3PkR
UAQfMAdDonWEnap6h/EzM9jMecbCgCCEDTE1ZYnRzUq7+S8QJeE8d1AHJZWboahw
TmGkiNdgoQW70gffTEzfVUq7eTGa1Cq2irYxHPadTHlK4BU/RGDYtKRz+UD0KJqm
hCe3lqsOInKC6I/Npgs6FkPROAznJIlVxSZORtlJpvuRQxR5aSFovLWAhV1LQIwL
d7w16U+5jP6SH54ko4nbY2h1a7gNnv5QaGaSfE80EgQ3D6H62Ul6+aXv9Jn4GCKm
tlIH/VhpmK7lhRVr2+k4/MnpRKxu0r5eBjtLTtCdeRzC6kY6hFFtOiJr/FFVnfJK
kvGoojMMmX1F7tuAiyZmCi8E6vyIW2iJpGqsLhE08JobZks8GbcS3CXcWqqLsuaa
5W3UCjpAmBGG+WQzZz0fcxA5YeF7u6CAduNAgumkQnrD1XZrvYdcQPEvOJfcdtPR
gThMfxaY7x4McK6+JdDdIBp9O8eR9bi0xfuXjWvAmEndxY9EVN9CNUMJ9p5epYBf
yVEBgyFIe/RcUXok7aqjlFilBDvb6FKJSnoWUxAfSVfWP+iaDmWYz5jLHsxPhUwt
rTxNPeOZG8GQl2Bft/YgM0mfuUhGci/3sfEyZCS0jL3x+A5mj0ygOJ5uuyzL102o
shMH1aXX76i4vAXLQx7zZibME6lcfP9C84oVYSi+eS7lOSaO5rHofc2wdX4WxnKu
xBp3ZKDfrqKeaRc1QMK3ZRIR1iRBI5jZzF9R1VOo3nd971fyQl0QLWJ+LtYmjU4a
xDCLMBFLuKicRH+iOP7Za1KlIMYbVNPHqV2lopTBDA80LJYAxRtJt9cWz0zWIer8
oJwvSxDWKwjmy7sjTVp6vW47sJLQaOu3rbEODNf8z0Gnc7+Feyh4OoGbk4gAO+KQ
9Ky/qtjYjzQK61UJG3jAfP/6juML+8xgOd0PQENpVZyJmNMUMw2OOOb7vBYBNhrC
rky5RIMwi1kAxO+yr+nI/VGVH+tPfLC9OHa0KLitUamE3akrpI482AyJIS3mmxhE
dAdEvnfwRXoKPjiDaA4lnbyayjCAFK2Dje7E9MGoJHZXw23pP1LtPlooojT+JNuY
nOFfiRWQk9+ljtTOvjSfErAKHGiAH9n1EX8iMLWO156X1fFa5OQsdpemYtrc9DRD
bKH9oGfhacaWRsHcOKku2Vw3fByBtll+Vl3IZbXVPl2ejyUPN58AQR2pnQNY1BRF
R8YzB99CyIZr84EEhZf9JnzjvOgFbrw3NHlkQIDsCSmui5Pfx6tQ+OPMtqaxZEO0
IqkA6C3soJHR7w5SE2linvZzIHyqnvlSEI1U1jptKr7LQIDj7JvoJ3QC9zwnIdFi
ByIeqs2krOSOWtH3comZ3yCxNpu2OuUDRwiN/zMdU7fIZhLCQxBTRcWsgSq2FiZb
BMP+/P2O6/8M+10LqvRL+k0xeI+TLVLA3GsL9mVJopsDMvcu0yPMzuvS3xhFip8K
Q12593IH1si4MOBuS1yF8IYd8dOOcKTHZ1jKSQX2wstpNlkgiMLl0q1/XLxRtHmP
snoW+p34SHZm5a/uUBamtr2uMc1la1p2doI7xx7HvMRGb2awpvrGOptUqs1Y5J0f
f0zVinGDqQ/qdoe2iOIu2bB7nFi/GNesvKBqD5fyJeU3fmUnwIzFzP4sxxk6dZX7
jTEdgXY1artpzQb5P5J7PzVVIg1APrEvBz6Be1DRh53glGkVx2EGxLq/trvIJrPY
JobWjgJjz6YJbAjiJhoayUpoI7y/CXgox4cjY4reDJ27Xr5QveIfZ2PuvSJ0OotJ
EMdgdPgyrEYD3J97ahh+eVqEgV7eMhhgUhIPUohrtlXagYKv2EqdUzUAk0qK8MhC
jEHfxPRTAuZYHFc6gAkLoyoMgQcy0RaQTUpi9hK6D4p0x+enwcsICZ7GIywYpNvD
nmfA7JSEaeo/IOucm22NJqHOM3vOFKX8+GcRyIVoUEzs+91ShMebp1+AjO4jG9lh
QYfS4Q5umTji+kmNZI7pk+nc7uy7mNf7fKwcRNV1yXlA9qbDUCKLjDwd8jRzJBMe
JE4mL8nICQ+BkSsdax4GlhsyyNrIH3t3ASjbJBNl0uRvP/Qx2xh3wbvE4KgkC1Ka
LqzmllnZXn3nmhC+U+b1qxxyLmlXSZ0Xf9jvv3fvSmiWGWOS6PuZLmnTc61qfvs+
f0rVF44P5J1D+z5Q93B1Ktv7CaE19qjvd0P5HPedFdzmxV5KJipTaT6BRLMJvjxO
rgTnliwMgn6lGAqcwzPQ3yG+b5VjK8upfRoS9mQzSczOI9jc4cass8nT5K6pdVTa
wmx3hWR6RgZzRbXTum76cOm+dzrYLXvMTpQZDOVLGsndu0W137bM/SY7fluSjEmy
2AxSfjXe9c61TRhKwMvPRpgTItb7pK3iUeBQUeXsYYIwBgvyiyRlSZxYXEFkqIj0
WD54pM6KHcBpMIv/wLEsqq0aCybqMOaKqGXiO7a2l6IHRRF44oN6CQXegAaKmCUA
eQGTXi7m9w6VgvfTZs/XnthItndI1Nr6apzyn5VszTM/BipO56Po9wsdzxOPAmiD
k+hm5bn+JPAtaXnlEftWrP7Zia0HV+unVWkg3eZsXBj+ffjz1ZN+5TF/o/goBSuE
sSscNT015W9gkgxi7XHZfV9xGpY+SKT/L+k/jcklQd167n/6OWVv3GSSm3pmMQEl
08Uq93jYQpNB329hrJic1r7BnCwOZXIhXJotb9hZR/CWP5n4BXNr+vlDpHbddgt7
WkWktf52+oe+swW/xgga3JXbyZ1OaiRNcmJr4Buq81bRCUucf0BPaX4zuZ5epk4J
c+T3plw2YLg6RoIT8Z++941NYNmotk2wLdQ5BXBeBlXeqA2wZ+pkKqk5vbeS4Kh1
StC1zOowa5J4dIfYom2mxQtNhgIfIwu8PMQNi7gKuprFfCWaO4cRfMTObwTu37KY
tSZxrOd0QWYE8B9HWd4e2FaH1wgWnprnUXAJoFn2F/gB/mZ7Tlu1R6HNyDZRigHw
MHxp7N7ZoVCTlHCm6QltWb+j8qO5KPohKeJ6bvDrLvT7T1ywy+wx+NWNbPDl64C5
Ncf5akU0+lY3awkIYCE034R9jwQnuJbKbJw+kN+oa0cTuVUK9akrO4TNW6HQig6q
WjJd3m8BLuT6l14jpRmM0hAFS62uqCXiYKHePm8JofG9ewh4NyOh9eEKEaGOJOAD
ZJvdoFBhxzAxZDm4SWjchvv1ZtWMCFN/lfkLagI44sW1FdCYsburK5oMLt5r8dr0
xf33QbObauTcotEYJpigIIG5JTfXZsJ4thq/kp9e+YPbTG/dtUn/tsnpxJZwPMpC
gNZob6KjnI0D3CHSf9t0q8uuCaGdl8xch4Z8M4mp3GH36n6Pwjrt4dv2NKF1jGF/
eqmQiBATtRByPCSM+8sG2PGW9+WOSaTiDoE17RX1/FaAy0t/QnWyRPqhJhKfIT0F
SjzjuerGMn3ehyaH39//cGmgzLhSwk26VMC2HJNcKDnxgBqByvVeZgJmNstV/9jP
MXf44wsqlZwMV9lH3evQtZJg+ddI+VvVW66iFhaHeqgHJme7o20Y+QtrMNaXpr/b
WGwmu8BffSKiySfxysIV94n9tQWfVTcr9QLkHXigmR94OKLOFe9jYfSMCj4jor7l
WchkLFcDZ65+qoPeSKpDKIv/ni373qrq85Il3o9MTUi3G6rbmsBzbXAiEBEqM4Uz
ebYmOWbLrJmtyJnr3JVhstNpJTpOwcgiM6MdeS6+mrhNU9VrgGLgSCjcd7t7u3ZR
X3fkfmWCsAT/WsvurktQR/w/mtkJAcTCwDkJchacesPkwddPfZRwaB/L/8+Q8ctY
Zde0DsyK62K7+emWjAxB9deex3t0xhIP6UW3DN0rEeC1xzqiCP1tNfENe5PgJWY3
DydsvNiQfj1xN0jNyoOLuvhdaIoJlI8Qj5RlHDtLDPBSxMzIWVho+9hon5T8iFaU
EoANHo11OMng44kKF/KriUDF3IBQcdygzvXDdm2aveavcHP7LLLwPEDgC3ALvyfw
ZVLsBWBZLLKll4oOhJc3U02Cy9owfpPjJCOGomhe7g1barRh2MJzo8QlSFiL+dja
DWMQOJRFUDgWzosDqmU9f0AwdIybCpKxg0jpuqDOfhrDXO9GDgGu3rUapIN0lwcF
qg/b53YLcKbH6CS5//XgczWcgu9DyFZAsWM7GuhO5107gnmt8yIh/p7IMn4nv7yJ
WTHGJfFt4AqCHWJlZ51qq9YqYW6lqBcFcGhmmkNojTUgQlugjF+iwnCqo5715vaI
RdcG1evA3bM/E+fsda8gt+hAoKDS+XXEhuLGtwmc/0sXPVDoQO7aEIo1Wz1bAo55
9j9jktkMNdj6YYgfZ1Epm45JB9fL84syer36q5NjB7htJXCF7qC45IidCqTnj+Z4
uIh4+ZqarFqKzmB0GbHDEpUsc3PlfVx9MqFJD8e7yTc+/86NNJvyvR77uEHwRn9J
L9jmEQsNzA02KGtzDwOtFrSsiuESGNA1PwIu9sSGbmnC367u+r2OFwyvZt4vDFmJ
0fNSpI/4M6MAViw5jTq37Rs8oHVZRJmZXvpsChVUjO1/41P02dgbxSdaMbu+O3i2
t6sMQ+rUDllwah1ov9fRQOebZllTIWO7rfhTXNLBM+1xcD+kY9nefd0y7f6TcZBS
La9p3DQKMNL3Yq2gVGZ0dDuP+YrNJ3ypC8maoOq7JFvFpx7UYl3pIctO3cHcct/l
GpoN52yFW0Dq94sQERxpIj+Q5Y6azLyKbmjTyHzJa/Shti/zzAoJxzN36WkGVtar
G1sKbL3dr6GJeAwZO/D4TLjA4HJsd/ezqvU5w7TPqlr7kzqsBJ6iRL7zOaUWKTxs
4XiMxhBH1baSOQ8mHUoR/hHYvwxRbvd9vgi0bbekvbD4qUMNuRNl2WJdwq+4axPL
w8AltJvucryHqnmxIkWf1AMsHdlmSBUSwBtrrWWPe0W/JmgxSC3BUHpm2LsmbKIZ
emm39R/hyIPSFsz2TnUG4tzBSRef8U7DUrU+0BNBlHdnkrJSZJRWGzgvMNVV5IFD
9nVLYqEe2LEeyPCbXT51wnI+TjB1i4TkJsKahiPB3+tb6LXeL0XCgPwNtDNuU5w3
sT/b2lpy04iUKsjplb4Y73B8oVzsLfFIAsW9ntjIfek6XXBwdm/BOK4+T4KDNbJb
fE6eCINk3M9Jfz5HuJW/D0L4Dhy3p+itS1eXosc/NIQUnTVaLkmzyNkDKr7yndVt
D/duwIarwQYr8WzXnu4wsF8EpJg7TXz+o7aZfk4ab6a4UlL9ZNraMzfcg3mJwlAM
Ar9Wb4713os/O1Obg7NzEl54Yw5ls8pHWF8ojHQ5yaRNStWdCz4kiD2YSoJMSGni
ZSGa35+m3fOQTgqoRv2WeUr8pxfq2ELuFHHvRGZQY2bB6J4kFgHLyjxj0zyCKw2U
QOzJ6bNAtDwpCbndz5i8Swo+ECO+Qcvw31x/ZhV7O3rRnobgWXUG9rIRzGRelm2p
czs4MWJMm1GZ+i8nfewCskhKGTrDWIDQdy5fTvBqMZoK6gGbWk9ghfXkOP5GnUUQ
lCLDMDWUVppZuf4ctkdNcRxt4CwhQWXJwWYAy1Ugrhk3JjXMFDK+fsCPPMN6ZZlv
wMZU9AV9Tq99iMlmrrQ8KhkTNjN6lUX4jLrxSyCtW993jZLS/GxRjhYezm5lbi5u
chdidboLeHIXAnE7IllNeHlNWyLiYDg+HR2vBeBD9j++AIB6OCT+CIDJ8ANTx+PK
ADf7R5Gs6NCHYDz/U51AO8LloEJkqYL2IXKSpPLHZoRdCyYWQdZhDAdBxoS0cOyK
XceWvCPilDIxX7uGX/620SG6/xQE6Nx+TEsW+7Wb2g1H22Zd55ElDCIoIwbwW/CL
+dTgVQZ8/eMVN8Sm1edtpBjZnP7EAr/NXo0q1b5YnsPBLGL95hD8w8LIrf4wf6Eh
0Fos35WhDBldmjr/1hX2yp1S75cGS+IfOmg5t/86lJRXo1joC0D198RbqU+cQI2a
I+94lGoh4z4XQJCygyrFau7DTblaTa4tX0bbD5XXT5gUQ2AllwbUtt8dsbiIuQvo
IxhcAS1AK5a0xK84TT0IFXdvMfIfJcGJt1lK0Z47qIEtepRKpaTNCu9q7PPPVOrA
/jBm81ETaZBUMmG9+2hH0ZXJ+Q6VZGqpsg/g9Xa97Yze48Flhit7uPdGVx6LnAlj
f+uLQ2otyT2LmelVLtWkkmrjJ+8/PbgiRv2jRmEFfzq+Vf1aP4X/qE75y4rzpcGq
kSKp5uAF3zcjV83VIa9N8ypN4PhPzOqm5oxZTqg3Ovnlp28NyPMCOU26qIPn9s+J
Xg3QX7jpUEuu48/OoD2OURBWDfwWChRlAl2QDluv7FK4vM5N9hhiC0ro31Vt5Mr5
ip8qz/S+a9KZemB5afmjoqI6J+exuKxK/9qvWTQzyOI2/1Dw4Gn6twPVbkVW07ik
VrBOymNNp75eEpDDaHUa6l5/M4CzL6HErTStqJ0mJXjSS1aaOVpo3eEYBUwc1HRu
uxHELYG4XndkWVvzOQnqOJxEiBOc9i5GEJFILm8KJ6G+jLvDF4AvTsBGLxy+VbCR
IotDKfvfC6uLNbXox+1/Z61iy2OVvMK4Dy48ifp57DZQxcsq/b6aAWBIXYJvnjvS
VwZbQZ/SbLti0P7jTYR5QJAHa0qSxsPu+xSryQv+uc4dny+Lw2h80D+NXqhSHM/n
45BiRGsPxiqkecyrgoTvrNMsoxTfrd4ubMhoySoET1PEGLxcLijHlHBheQngcohR
xhT1SoKj42Au/lDHK9DRPrZUL2ikbBMeCUEmK9uxb0KOaLJbLgFOUiNoeCGQ2dhU
yo295CfiAwBEEfInsTDOgIOcQ76zeXk0Lwi5G6+/t4AbEHrT+Lv6ZrkKDWxY+eL2
olEDf737dW1V70MuyzG7ZTuIfTNT0yHDpDOwBmlQvV0L5zdrpFL/I/h8LKB3rmBd
ngH3UdjDOBvBRQiP96KQbg3VF57YZGBkALLgF1sGOC/hdTfYzCusgasWDQqYoPQc
WOmQs+xGUN2iRPRzboLHFuvDqlVNX8ldcdBvEhFbwaAdYPEjWck3supjQjTqhlmS
c2Zc2P4izEWfytk9h4qLc2URu3Gmy3bjniLrRqX3fb32guS3kJq0xHmNZY6Fh+Fo
NqWVT8rGxA6VAeMeBJYX9+KVIZI1L9FrfXnQO88IFKHZRQS3jy2idu8G1MS5typg
LjYRoiVbwU4mseh44T22oKMrtmXECyV5pimfM+vQNj6qi41cWJRICYi+cFi5njjk
p8V2CYlcVSjKv0gzaTm9iBV7lpvCgz6bqphO+1MK/tZsrHRhMcOuv3tv3Nla+S8Q
aHxC7T/NglMfttZfroBoEoQluKFZwwNTHNF1Pv/5qU2ePVYAy77b9HmtYb2cFD0k
aKwvpTc9QOX5oOBXC/yxZKZUevq/hMP+fWyZU+T9WQFeZs2ZVt5i7AOLP4qZlpud
LpGSCRpDNtaKFX5YvgV81cUDamhBVCe0GGNK6nbzpa0HW2ou3x7b3FlS8A6zrQJD
YzM0kV78VvMXqM+rUpyHJgeAHdEgQIZIByJxnwFOCVKyTD1f1YtoprcRGQ0C7EQj
SrU4Z/kpjz4XHVvfATlRZ9YtzeOUIbUS+yHKhbFQM1r+Qto1/m8UpugH/oUA0r6W
hSx1Pv1agD7lVrU6vKjpsr+hqtRo0fhqpqr/0DlCrmZ7vix1oxaAv6YComyvWTEP
JQ+/3MArR06/vfZDbnaImB2l4F2rpmvEuO91cOEFaYQIpha+GtFZCKTI/f/PU1ou
kPh1gAK75cjtOsQAx+Q+Dr4TK/jlxeO6I4x/EAy4N2NCUw/GQD1zs2aALbxHkXJo
H3NMekYQLq7wfoZluz6NwDl/lIixfrs/zRETwQYvlLCaao+djflStu3/anu78hTU
PbLrUEQuyHvWwJ/ZElHqvE8JJNGljgZUPiIzkZCfvK0vIy/Ox54xGEb5LIH/P/yr
dNKEJRv/PigwdyS6KsQAhLeojlmukyb3n09AEZVvqtf3QqEH7jruZmfEe/0PQ/5h
MzMagL9t5orHNi1NWKv/RU6RfwKsOtWYvNQ/DPkFUPudQCKJqjRXYaHHp9fDoSqr
YMpinkLljLk91+Z92PRy/oeNIO+vLiFbtP/QsOb4al3w535CUVPZY++QxsRC+0oq
MqRRQIEb/YwxCAM/ZgTGwYH48CrBns033X3L6ei1Q0fYPqCsTdBHxjd/6mppVIiZ
JvJti3XN2TM7v4THwMwfnHGR6nF3yzP8OzAWLqUBzHcX/a0lCg989aD0GGI08sjN
irs1PauU7Mn5J2Lwr3MvCmhWfxhlmBUOUsmkylb5rIyVAtNkpFQDOlvWj9eIxnvw
DtIa6op2bP05KHP7OqoSJGWK9WOxGzUGygZZ46+CKNfN6MaMSSJlEg3M61RXahbU
2FluuYAf4t22f+a7M51w4Qu4945SaHJdZyZ4UGep8JsWXb5Bkqdv7I2npNpJDmxu
tS+RtMW36fRs34n7sHCuFLQdQmQu5rMszc8bw4XPMeqEJwS6THdKkwmyjKPHzNQT
Iw5/QA642dK/YBbQogTnU0QTHwV+T7tjF3eLJ/r0b0ZvfRLfPUQwlfoyEfjlHCjT
JLKV6huUOFe4tDkOGGKPn8xj30L4JAg8BPncVqkZQlqo0/+oOiPt1cH17DFcNVSw
tt/Z9v2CPaSO4brFNkC9ZGZAPzcVJD3Sd+FDp1nZJ45hizawjEoiDRafu65YdVwO
qy2JX9wnqg4rnz2zh5fD+kPo/gKmb97SlPVYxTC8YvyRXJUXe/inoxsmIbivzMXA
JNSpWbR1V7D7+K4vJJoask4/ZyqzCoIUK31tym2Yk9a75KPo6XhthT+Hm0zi0Z6f
RqVwWDmA9ZhWgTH8JmT/VagX9prQo9uIQ5wMv5/jVpByrCqeUn6lN5I6hs1S47jB
FSbNCcO+/WkUFa0OM5KnsnoVF047ZH2ZDXRKQTTXJRxwYZOocLebEa0tF2uGcRE5
S+0YsBRKiJ/Prs0d1e/L4TqSehe+YVWgorhsQuLRr+iWt9HlZF0CYaHBG5x1NyC/
fqwiZ+Q8Sj7ko/ciAHoKW+T1MS+Ia9+7aU7PkoLW4UauQ3xLZlm/dlifaAjR3Q5j
JQEf4tehQngZ62JlEoNuiS7nSZA++o5P199hhDBVYCqXfKRdDg/w5w/bzbTRoMq/
`protect end_protected