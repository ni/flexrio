`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 24224 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
YachDS4bpHRDzLXFQC4CtbQ03w6X0EfT2NdpchTmfNkI2MretxmfRNeWpNhzN9hn
XCqo21lG9AN8u3f0LQDEpibOtQeqr0qQtkslHhr78MqZcvgJHgHHGj0628PacZl1
ooBb24NuD3b+IjxQv7xN3BgmyAvX23y0ZBC1ldrurTUljIWJtSy6RVmZDvSzSVrn
uzqsJDJ0SYqVkrvpaH0WHx7DfsgGS04g0ayfJ5HOL6TWDhCdv4sFQeVA4qMltcrk
aGx9ksY1SFm1vTZvwtYewdXTa38Fek1ga9Eram3J/HkH08RCAomeWj82mOjB+X2/
AN/i5TWrtdtElEZst/NVb1FTot/1rdv/VvbLpXK9zVeadWvHrIOAA+0zTgQr8c9T
I6iQ4D4cXfkuOWIkiHRdEhwnclAJwQxvYjQmoBr2cDdW4UvZl+usZ8BDYkOGrmNC
uA9/WEJrVaezAY+dV6ldJljJGqTUf69WUFpKKAcT4hxheFHcKsjNlVnePDvobZYI
RM0bWBJoJZcoqUOTLfpNp9dXpED+OW7Bf4nXdqhWghch5bqhNxVX/zJTTcKPX/LO
LGiBSYn5cwwvGVPnhhBeEDCGZiWwn3sbGu56n7NpIec6bk2uOdYWhzsUX7DrEkgu
52y66fWPr+I1NyGl1LF1Nh5Hs5h14qWLmOTTUY6Qz1QeJUf4BP2XYTIIEbTjYeo7
Ll47XPjpqTnfbaS0atk5xgtS8gfWsGjMpvSt3GaeY+FpZDwmGAzKh8oYZAhtAYG7
dBeI+uc7MzEArJzgDY1Td0nYwRPMRpuO5xJLJiQlMcglAfqpek6LjsfbLc3QVyep
nCxFovfvpwqSi1hgUvCMQRTHMoCKQF8h61cUuWnUlc4UQq+JTvZAck5VetSknQKD
wD8d7WzRMGUe6nyvXf5FklUqrhGrAdSJKfrL7b5k1VoJtaIh+5mHC0tbKdYODd1Q
R6j5LIdUJtop2E55pnIghKAfhDrf4vY0UGtcVR5KWGRTScGGTlSQ2rjZ89vTDXNc
DtFc8qRE9dwDFW6XP4EQGzHURCG8OXphR6+YV1PvskKX73Oy/3YDrrXLcPEkmMJC
CbSQIfsUYXHcWlfnNJeKzcIyg1TnS7jnnxGz61+4QO3Ku2FWcUkjmkDMxGuBqlXf
/fw0P8CpVGCD7GbL7qmZuuE3VFfX8QenBnLH9xC2Ivpf4H3XHKhTlhOxOQALCvLR
N2QujPisI3I+fXNnjbLXcoM0YKjZSFD9UwdO00iUH2wMhJIbwJ/uH+e8HJfovwnq
OJTSeNndrsdzYoahy/Ionxz2Gfx11qVkPcvT5qzpcNlGOZeZmtzsKfynVGs5jYvX
W0En2m2OtNqRkv/NU/d1m1bQD9UTSgVR5uSdbBptZMMU6kWDMPbuFBV2odL4EwsT
q0phz1MtVKXb33O9f8m/CXJmgAmQq76L06bRxfstu09vOMfD3kBojQ912gdt0JZB
zIltG3un/imBq5zHxflxgxkC659VzEep7pRAZZi1BgJZ63sLr8PLO0qLEH5doy1o
qvtAYfD3SKFruf/M2ZJu2oJgB6RmlK1PA2LuRGcEosuOd3QX6cSQ5lhyVzgnb0+8
B2pp199T6rtTG137+PWgGGx8e/kkCfHWdOczXZlAbEntGX/fdjITGBIjFLGeMyhI
dN4ZHboj/67WkOqdddtjdAzGLi/c/UDiD8HCnzlEMWOrulJa8DXCiAQy9H8sxSdY
NoaCZlN4pWxeNsQTUwihzufpjmnGPx0S6QwOJqhnOYXPLKSjxLZz53yP4xxftDbS
ffvHQNIR082mB400scYez+uutML03rgJPA0WmlGyjEXSqeDtiCNFRykXzxXfz/vC
vgGJJsrLGU44iBnMi4zXmfD4/zRbeUutr4DYz550ubhtXkjs14bZFONmYUPeFsUo
0J6EQnNBFMxhwMRgOzFFaWNG78epy/Z1lOK6BuqxL0+Fkb/H+q1uXLCMGrnVWe7c
BSRtc38tpR9Cmes9GeF44tJi6lJJdHkPRDEtcugvMibzpOfa+vfWvwnnZrRqjsL3
drxDRCskQ5wCRoPRVs1Hl2cmrD2MI/p5QjhRHhQM0JPdcVTqxCtwmbST8BT3o2El
KWRafaJPhfUu4rTICxRi0oW0+ZVEm0r+/lst7ze8LU10+esFtZK2Ze7FMUzGkdB6
Xmtz1Du/T949FW+YRwfJAFRxB9+Is3xTXN+z3Z14qw9ZDjJWNLU9LeHvB319uqUY
p2yb20wD3/Ak4xXi99AtI4F2fnj31SE7Y16iDx7NXCoT5kfAO1S79RGbmRCVp2y/
f2oMhARHox5kjtY4TWrLAZtPK+ZSwXDAwySA7uN+Pn/BqgTix3HU0Ai/PJVl+oOZ
zWLzoxqidi86TBPlAS/DR2sho/MeshV6vwH3IPrURPpfMBdmgcKAk5G42zn5CQS+
yGC2hdvz7UlMaxnKXwmN5LlVnsRfiydYEz/s83KLDOHwWdkBtgohyglkswdwgI8k
/xNZMCmTmr+s73GW4tDHCsMFM+sfTcBO/Vd5OtAEloQrKjzrsqN82v1U5B3bH/Qn
I8uCNTYIpf8ACeAsHmhnPBwuJTap/LpPNDErZAH7J+9F87ZbCfshY7IbRdYJlZX7
qH+YGyNAk1jStRznSX1irv04IuC2EBVM8+G6NMIxAZghs86YEC9gqnGj1j8l6OCA
F853mdIHv32jp5IaKNluLkXRwplax72biNNvr78NKRjg4+VGSMsHttAI3u0me3sR
Ufa86KXFnLunfaq5TYNWZnevw15RuYqHl+Nrr2sQlGT7FaHkZyjC4V+uwjZH8ncc
zEpkSK6t+9r33z1CwM+vrCCcfPq12Dbgq7Dua4FsvYq7NQCaT/MsL6fG/1TdFEF9
IV2xM2ZS7umbp6vdhK0OUtIn/cqz8pcJREia4RAmzY1W4QKGOOFgKUZsv+1rPEDm
MHEEhF2WGn7bDnE+PUcTHBHOjiurGAu5Xjpw59hDqe5LWXu6tD7+mpfC88D++N4c
Pdb6/hHg7xv/5m57XNd6Z31eWghJ2Ss0xCzBPIdy54WNW96itQL2XhBUDrwXyYl4
6xCH5tEMk7Rnfdpqnfhyu6vmFe9RUbZUESnBi8+zoc3gB8MVtzSUnHoy5SFxJIjY
Bug7AFbIbxEaXu5l9bLn5ml+9tdl/fQ7n1JU6vHnfgsvPiIXvcWomqSzuNkz3DnX
wIL4oIU+NDfutqVG9tANgpc1NU0F8h8xU7Y2ouHIjv//I2+M1rN/njwyULCYnZqE
Xzd1sR8LtTCabq4M1VgGr4V6N97v9HhL4K6aj+3m22zrYWZkbO0IjsbvmwMV8T3N
1B3UnD+aU7ypciZWiyxtmFAlTqSshJW+BcQqbAjaQHv07dGWO/ijX3ecDU/NDhwS
MAhDdgPaXGWRy7pp15vEz+J3dqUai8P4ga2G77iWZ+UwMdESsFxbaqBTN45JYKBL
EJcu+zhDeo2Sz6mbj+Er1HJ9cAsw+DRrIlY+0SIZb8L7uISGB2zTB5D4XM4RUPBm
gju6OOiUH+NETRl2R6tLuAIn1C2KrPCEBLF8V3zFowZfbTF8wP4gpOYE49PzRnTs
lxbYjqnow5yQmG+g8nZF4aWByaOXkBo+QP5jfS73/PuhHm1nBjQc85NwrYBM85M0
HhvzUNNDqlbugp0n6dTncjguBJe6edCS2PtuCYUQS42Nac4cI3zJLZQWrlPh8mK+
hDBpA/DkpdNN4OIzYPj95K+ok6FzZkh78Crdp2Y5rlHysjXlLVF0PSPdEjUBP49W
+p4DtRtSnUoJTfrxYZj7giT55P4JOVmjMBN1OQe1/evv7+HWlmtre9L1GQfw5SJE
3QgQU+3KWI2HILbHO0FkiQWu8gO+4RC+qxpeh9dt0tlvxm/Hdx1ZXbQVhNEwLPS6
nfQZKqcKsIm1QauoW6mlaV/eJnJhV0bWZK7J/t3VqtZoizaYCswqNhR++Ye3wv5u
oP5J4n24F9AjXGCGzEk3nSBMZyjcXG346UFAsxiLEuvzZU0mJ2+/7ddsDpr9QJBm
XoZJ7oWqWc0Wd0GaEhm0i8b6z6+YwcKA+9XC9buvRoOsHd7ayAU/rKCRTBDNNX9d
wZBcd5cdBbJIMeu21cprtf7A3GsVZiP517V4mcX9L54NeyKQ1+LDhQP8tfy2wcRT
D5Y+KOgIsY7OWgm5Dx4NUun7MQUIa6uxtCZ9M7ynOGt78cmVmoe0Ww4kyb2l8XhR
1s5RPcqtVxfzxWm8MGRalgG/hFQyktx6EHUshsLJtCieWp1WqVJmzNNaUkLi2oKz
xcjK+fagUeAGmQavEs4HEKQAsLFE5ZDcP7NSgu1bNYNfm54izUg2UeHoZWdvW9on
t9JLLwmqjoHgcHRkRKPu84aSczf1xVVkyBu6a51i65bZuM2XbN0DFNpVodQJ2uWj
4BuIWA4V1xQsdQavGDJ5nubBgGLoqx+lQgAQgkRgS4Pp1vbjF7qRsRUWOehLnyjb
Zj7wBcC6Cm+ET9xZ6sptQhmIfAVCwBz8yVXPtGN9FZaoWvLhl4oY3ZnzLz16z+Mb
qSsAyPGb1TjygD5jFq9dmIP0KCWPmURUVlt3ZMVMFS2rN1nGxuq4Vanm1pdwMT9S
BUlxUSZgDJvGX2ZInQicNVuMQ8vtu2PgjD0W5+9ADhzGX6WBUV17M9zfrzzoQbaL
h3TNyXfoGQsy1dRbmBK99GG73o0pjeZRIkfzHEJ8dCGZkXJI+WqQIXwJ7m7FAlAc
HMifeA1ZUOsKTJaWE5jjE0sBHxjjZqfFnrUvElWkpqkOYZSS5XoqMTmYXG+VzZpb
z2WcPgmyZBsY9XGFNsmjXFiOuNR+/ZtrN/bnjOlCLHnXArR2BbS6fCLAik+pAkl7
/TkVkzvHS9OO6471iv9fqpuH775ie2Sk9EgDzbn9M1uKrpJYaU8I09Dc+tOWqWl+
nz4pVLlnPZuAeAFsFc9/pomvK528b2CuOmKQ26s1u8bEvl3sk95ah2xy8FLvkF+T
xFr32lij1/pBCNVQ7TYdXX+U6qA7i+HKMrnAMcZUB9x206AFcb+pcH0uhjKN/w+g
ip5aVqqGfuDDCQG8RStX23OTVqLalbAURNMoCArEJdL8Pr5FyA/unEr7Ch/hSYbx
WykuSjuTkIuh6D7N9voPXxMUjmMgEM2KfSMvHBFVKTzjzztVpDkm7aO08ju3Zx3h
PxDKRVkcs1XP+/yYVZXPVp4HYnm/1TJSuLaw/v2m8ctFNJTpIKYdG14C1wDvbPDh
iOYlbnGu9F5huBTkMvdipZMQfPGQunbtZU+Jp7XE9UJTHACBfFsZNVwaT0Sf3FMQ
2euOiTVq04aW9KX4FKQz/s1a/DAU3A6sDtMfHeR0d49bpLvWveONNY+9evnbdwHI
aclJMeDdeG6aVY4iMAC+GlIZnpC87c/rdsrB8EfPmha7HOHIwH0FLMjd2rKw0oqg
stH2iZjZYBQ67ukPlVk2aRwXAhq3xSf1VSnrVKSNL8GnC7oBU44l8FhPh7FG/XXj
UtFl9SQ6eiqLVGAfQ+ep8mpnBDsPJizhEUVI1q32xaJmnxc0UTdapcDPHGzVgHHB
GRugnytjkvIEHLfAoIcU2foBfSiOpLwfaq8zbXeKL8PTP5enY0Afrro13byS1nCw
WWpBSga4xKE4KOD8MiT/qivpu7unuJtKDrsw170222AmVDgxBKBRhFJNo3d/gLN8
u2RdsUXP3kQbVKkEVSo+c/+EPPn0acv6ySXfcEnzpU7gCxaZDT9JlCCDh6hM2+hc
GIwABmNDzEK+0yl+G1NlxjqaoFWpDEgHzcDeO1IoR6aBQQBpnn21OiOYHTVEBGLS
HeFC1BeKvIBU1SyfRxC+3KEuqP7daWWOPEGznW57FhFYP98BEg+5z3hTIsO2auKY
BREgl9Pj7tFTtMahkjKB/as0M4QTOJ+uP80oAnyqSt3/7hS9upEMlcg2VUlJ8fup
EQsVUhXw7VwyNpuMmzPXfD7Bmb6A2jgToLMvddO/5x3ed7fdFyHx0eFhGQcWfkdy
bXdmMyBZrffgA9DmRSuUswLrVfhN5EdcPgzujtJ46g1liEf8gChRvxtF0t7C0GCW
QctZjJtGTHIYBrGkuvDBoRQAy2/H2mFVBTTwej3sp0Ow2aYImlS/RIEIVCGVRGD9
vku8wp0RlGkoWQ5zPgoObmotA7Lg1KEDg8WlHv/OEWLVDt5zMsy+SOmzhmftrZCe
M8jtX2bd+m3fDFTLCu+Ipr45p4cYSBIP/G+6IYcgbZyFx4nEnwaAGNu3gEB35w/b
bq8p6/07Fi6ZLMmeQxXpUPONKNX9AeuX7bvRtV3G8VxdElbAtEp4WDAW5w2Tq4Dx
zHQC7gMlNWUkBxRgAFuUwjdjrCtkDmGdDk3asWlJwaXm0YPaSeKF33iiHXNTzD5v
JNmltIystPiVcO7lVOkT3meauCJmshpAuO4IqictbVwp1XsFRj4fAqjKXwQQzSOn
yPaYsByaz88T32GX6Ynp6iIUILqP/Z5wdpyMAXjM/F3bkNdFMFs8mIAqaxQOwnJ3
zEdAN4bxDOusZovRInFzglbczouxTLDYoLW4LiEr4vnf0s2lGnRbfUEVM+4bYIZ7
86dcv8T9I41BBJoznVWUNrwJ7pFE0T1Kcu8CwE8lOocjxvqbD2Fcmuni3bja4Fd4
2wE73UIHcYB0vi2ZoVsIV3vyzNXwF8wOZYeur7kqABrJpIpt7hLFOpPemOvs+YwO
w0Zselu8S7V2slDaxULpCeX42WrWL7qYvrnNT137QoCRGV4snT1BxtaY461V+aQb
Ce1ZmTvJ2JVLo5XMFabZpFxFAQRbfgkIE0nWj9q+VujY61Wr13GuX2ZVOnfLBAuz
DIBJHVPrWLYFEpeteveWtRQEpX1StYODie+lKFhpfRhD0FS7jIOggyDmEAvPg2d2
j7AF7jWJtcTljMMyIvefL3/B7voNAgPD8Mr7MivTbVZvG/7jr4UVe515OrYO0rop
+9y0F4uW3fSUEACxeZXSTPU0qI/lK4BeiVb7Y1ycPpHKJUD5bk/bfb7nNaStV6eN
sPZ3AE5wFMgnDVTOYGyten/ysYw/KYBHKLhdtmJKL4IzOUucbKx4t8lkziQ7fTs8
o2m+BHWD4ouHIoAOcVHzRwsqaUrlhMAqsOpYwzCvnXaypopqE+gWavgxhdoPpFJr
ZZsv0o4PvV9QzOeSVYVxpaPEHXOr8k4IYmJEg4SGmtBfjYyfe9q8kIxO40n5m3Ib
Eja10iXhcXkSIjILgHwpk3oT+I4ua5IJ8uz/UyOoLQ8gnDARCLUTmzSLjhUWhajz
iIDWQbdd/cceG5FRlkxaqXc+vLoo6yS3FDQ0MPciK/KPtB/PNl3HPq1qR0WmNg6z
7UPRBpj3RD+sXhuFhLvEP0qLdxu3kRxrCRstghs5E7lof7Q5WKHuOIXR4I94cGNj
0sXYomuJCqa5bcW8BogPJ00mqc10QvqHLBXDpFUw2ZeWimdfOd5L+YjmRq6Cz8/R
GGgLUwUfUCWCtL1KEZf/rZrEFoPei90uNuqYvgViyKlwnZgh4ihuc9fG5ic66RdX
v13mvUgY6zD6MbzvDxhvPkt3UTne4TPob8Xe2KfOhpcPlQXbUcCcbhlzkHLq3Awk
lI68WJWwaYpZJBCIEHLW4JQ9AMOCqvLh1E0UzKOn++vH1DqvL5Tc4BhkRvw+rZXk
1QlGMWkK7Lliab3TMWmzLjocZsE/kO6dBGJncs67fNbSxTN+UeXKoya8Jg1MS6ZB
SG4OLh333cYaHjjlUu0ZQwjz0yCBh1jlBqgYPd7lY3LFJcgKPM4vfgtuSJqKMSc+
qzH6AgDayu7tysTIo8jAwkTSf6f6DrhaDWL8BZ8OG9KqFPqlysmfvAb7QQ5MOOhp
tNuAAL69yHlMSwi9fZ1mgCs3Sn9fyREFa4xkf1R/mVqsJZI9uKTR8kGOb9CAVVYx
AYAQQjtJ8KRIDHb2Wfzjtq1TGb5Nk99bULpCksMa1GeV+wWQEj70SyRCz5z6W8UU
U7mMl3Tqy6CAjsLXQkgjzzKrcxxRBg0XerzHJBFFTXvus2+nJZxEnrOHpl4//l9k
gcnZD1Nrk8XzA/6csFquRwh11lO22rxO0X7kWaqY46wc7jvh5V6vbFZMifNJYhGp
U8pFFv0U9BiAiUKnAuc1mtptlN+lfrN+C41kgg1ZWSzC2mwjUzdtxiB3J3orIC7a
1WHmyudU/sGMV/QOsqoomI17kjPJ89vhwr/myqSe+jEA4jaqLx6rhaJ7/EBTK4H9
WUXfedV6E3TIE2HpK4hz6dEbSTc4ywcho2UgSaghu7As1ArYEKzuUHAZ734OiQtU
iTLtdwBuZVZtmGVTrYv/srnh9a5LWIE9rhkl6Nb1j84fHHrbXRnRQp6jBGb0QSWN
Vu+yoRUioQ2SBrfW1WM48ygZt5CSlBcnjQz1DIznTMePHTMjSzGLFjK27R2DfwwA
CkNIc8UNa1wsuzPvqmxjHm8LUE7GCMM4EyyFbuWgZN/apNzzVPHdMjIi+zK/Bj++
a6TMNqn1G0Ghm4lcysUD2KCjsB6dNH5BePX3syUA2YThtSWvYQNfea5/owKjMWbQ
bMn7jTjk9e/vaw5zDGAu5JjJMUWrQjWn11J940+yjJSiwdFfpV/xSH+mCIzojWCE
EsSs4j6X15rIYOMX799bcFW2IAzT7WgeJIUntILIxBSUwBqoUk29+jfrc3wjO/2O
c4LyRGKO5sBuR5bNiHQSfh0c8Yw2XJ0+hfk4V+SyPi8eHYPB6nU6GpfwUtO6hPRl
zrF1JDpOP+o99LVlKu1ArHix4csgMxDp1wGGlOmEa6KTDJiKj2y6AhuFLDXZX4lP
EDMauYYN3E+xmc1fzAifW+oHl01YRnSmL68A09GLrAWRUYMarDwh9NQPvPua7No2
GuhDlfKTj3AXDYZE5FGCHC+4rYp8ftKargxHsXaftYa/ZbhAlam4xt95G1T5OXDW
Ou+nl49vcm6H4rh8foMRv6LKQLA0r0NSYMfIfxWkyxKxB7fJM3SpKNkZ3+F0fmUR
SVsqtMKK99FeINylUhL18pKMZg2iqNdXEyZu6S5HF0LY+MMEJZfH9iWm4uVzEn3A
eyoEPPIMcLy1pqmYgshgajauMxIzq8TmOBrdqP3RZOqSuMjkMYMnoX33hfx/Ahyc
QyFV3//7yRFL5hAfQ1BV7WS7wkIGLIConPLfp3VqlPdLJNFAjCFynrd4H6zHxtlA
X5omFGVQoS1zDu7wPz6IqYaDJ2GpMvWWLaks4WrjEj9KOLwrqWC5TvAKfSRPd5uz
+QelK9MBDBD3YUvhA5vbnyR5jBgTqkZVNfNheNf/t1m8uKHZ4LU9LB20aUPtVxtd
I5Hm+v06Om58ACSMWIRg+wgB3pi3RjRbmp3/etbE0jhrYgxtr5lcGZ5rBjfCVinx
1ir7e6tlYwTYCLsrlHZyf42Aq79Sk0wFThuOMra+UCuyoArjGmetM0e3UGpQ2Cn1
HgKzSkB9rocmvqU1wZmIX7Yn+o0E8o0lKDRpvA9fZJm5c1H8O1uAQm85EZCXwbuZ
6bo1AkKLq6YqmOX7adF8HwsNNMDLgDKMyPuZXP0SwWcNA2Owb0ubedFvrVUvXjxu
gp4pe4vMG1RzKge6/8dnfM4z4DDc78L9fxnHhhPBFelJL2+XmUTzlp2EdIFpg9NR
R7iSzaf2dIQkamlks+q8jh42I5Pl1dNY/xVNnVcGew1IKaZw4ivzP60Jv5bJHL6S
qWIXK2XEDKEeh1xcD1blpU7s22tGmnFEt0GMRAbiFTq/CRBf5t1aM/wpwcdHXr7D
y6/wEUuoFF/90rBXcc8guaDVZFARDPEuRZd6OpcG41g4PJUpRiRj7aV82PuBKLsT
8fsaeKFQwlZgb0McWFFfSF4KaxkhJMK7YgL4d5IXTx7pNJb2sOxDc3PtjfHeKsaK
EUfyRkiLi9LGYHdMCXmuCZRfKQGxx/MkKTCSGSE46sgOTtNwv9/5GInrQfaDDl9C
+OFOrnvBNrkfSiIkDQPwywoE2IXvsb0lVhgfhvZwXlGAJ/SesOWZTqtO7mB3hsuv
6PLZKwZFE702+UREPxh57nLARSvHYcRDjmFGsIpYoEs/0s+KaVkXrvprNBIxwHe+
5/A3/4yL/PO3N72tyRzExjkF+pV8HDbgW+Se0wv5xYTjIRWhKeTlL3mY6myeSZ0x
ux/SeCFe/a37L9LTvzdRyfPIOot69M9nFSp+iYEpTR3VqwLN6P7MDn5Rw37WGtMt
aaTcjK5HzGBUCXC4Yti/APP8SBrNGOWj9FM2HKjN9gHKEOrUyfD1aXdJMHbYpiWF
QYt72ckpuota4LKgKWz2I1PMixWoj0g8Efp+qTIS86PJ+jV/XlQSuvYgtKwx0nAf
QvXlthD+hLF0RnsSItN0dGW2qyGqrJJMeS7Hkq4wDqwk0pjGJW5cgWguHJIYJiWu
1i2Wzn3gMQWNFKVoC0glycT3cGEBiKOglnHIhVvK6kJvCsNCjDIipXO6rlKfDFvy
GbY90rET3mMdjA+/9sxidG+Xlw7N/A1JLnn4jM5L2m0E8+dpwgSUAMw7g0Wr7jck
zp59h4FUCNxPwyREvGLcHCtQZac5NQPn9yZrIgZYFQDwKbeogvyAP/p3QDPmdF2s
k6Nu/sILIiSX71MZMcgugjmmHWjVNaDjtPSGiq84G81crxszgT8t/d/xtXWwG98L
VZiXT85jRLsxZZNwguhuhxTj4rr/i7bGRi2xhEJX6vf/9+B1n1XhSP8NLLX+4ZKF
8moziCUrvqvPN/pJv8D6lceGjGVceDabjP78mKAG0xEHem0aq/qfFIznwcMo933a
Wo69OgcP88UlriUcsZC3YLShU0a9nHU1Yqf1CxwEMqhp/l4OZfr9Y3KhEtKn3wDj
AJEGrQGVD++chzNgjv1kXVUdeMu37uOnMy70F5WOVMyoBc51pVwRxI/2LPorjXij
wD4iH8TVCM+O6FkLatNpr7hYigCLB5qDlwEFrDozTeDpl80ddDDwMJY7G8lZrvKf
FV8irlOBxbUm/xW4gTbMfrcZZ189t90zfC+nV3fBz9W1Tbb109xSSZ7lP0myxODm
xaCw7IGMS43nHXRUqLZ7lEw27voP3aTs3EZ5vWsV+7xTU3XSPrOOrF+ielCu95H5
cX5b/T+9F3qRANpqDrsITfGSfTFLnrC6fEvqVj00994Z/WpwHYwDax1DnAGTRKz/
aEmXGSQcg36sfmb766tNOTA6bjYYHYa/IeXbMpUxNELQS9fAyjtFOfAEFMUUm6Yg
GKN8ePtB82uuVSFIexMzRKbuzrAxABdjGBfgiRQweiLI3RGfymYWd/v/rzebRrSd
LbmHcmcW8WEDdjQ0Yj6gDZhmgyL2YMh1QjVES/blkATKG7pygrZMC05PsgsXn7ou
9TMCEjte2OS8keMMf8RAeCcMlNBHlhrtie7djEZ5yGFZujAJMFJCIYYs2ehSF+lu
F/iQ/+ZK26mKU7yNpfjt/0ktmEwuWTNiCXL15PLuKkoiu8UEToM7QGYJQxwOttKI
I0i8EuLdWzgzcetCZGuGOoESs48fhNlIjpOmc/Cv/xSFv/JhCU/5UcyfSNQQeDep
ZhkjoCQYLTi6y5lbiuzlDdq2edmAJ0lxvrX6psb0J/lJHddFHrBB+ZvIeg23qsna
Xv5wo7tTMFOYvCj+RBPS6Lj7o5WRWcwWSK6A/aaILcMMDqrKG2jEAg13fRdc1Rp4
4WOhKo370+eXk8wjfud5puFwR097k6hwFgud1ToTvJyjqiz1knKxDSD8NQNpuER8
VhUjTIoIvbiFAM9Tblpd6IBLVCoBP8hCfig/bVrUMaQ7sU+O+o4O1ytDbpc0L96F
uKhrLgw1jSAxBtQh2xfWJ2j2lufVhhe47GsurlxUUlEuXUyrs5QWUukrI98xG4OB
0AlvsEty23DkyVTex2WcEn/EBIbC0URou1G50r2whpNXJf2GjD8mA1PQZYpghcZg
qeJl7U+OBIHgQNHa0rmzrnQWklFzMIaYhrwBFGUrYJ+c6oFkhNq+48Rh7iZ/zLm9
4E3dxOkrL9HTHM166i8CBjW28FAcBLfw1Rq+BiGdtLLpiZ4GCy3DU4y3vurlT4cC
kvaIdHfvAvA4z1uRPNiptdQn9G7FuM/Vav6yd+bKCXHfWrVVjXt4tIcMhKKx6wq1
dX3WwUpmjRe/ID3RbppwitCZPN6zrzsQ64Z/n2vsg6tjzIvVQpq9GUiF5uyJcmEA
4IoKoUUPYT/eMvMLCMVMb3ShifuKWahDmlCaYOkdNjZ6C5ybUCHHJKietFKcBpFU
SPAGPQivR8g+d0RRq6rB1K7XxRBVvRyb5PimCSOI8HVPlalrqUKtsJ19QfVjEzW7
fWfVv8C2DlkWdCbm2/us4wyX1R3O4zZndb1K4Wxbuws9opP2Q1ejgzV+ThUB0hIF
SztXo2QYfH7SnBWLGKaNHC5OWMOTKv2XtaQ8x8f2HY1r0nIe8Ek77nqXo0Bm6nO7
lRS67iQqeunFzUwmbM71ZBIoYUoV+sWh3+9p6f1I6o3qTCSMnKyhp25fB9HvubPG
c3NI/3aiUSl46lXQr1Og6M65fnKlOCXUdncwghqr9BCGTcSlT3Q+t6Pn6nwyjLlJ
tLt4kQC8QCbE2jslnpTlam8FtWuX6OQX4W9skcnVpWhlUfWDPDlf10Bm7ScYwq1D
Owgv0HovYZ2PFx2uroXGWxdNcM55jGGO7LKeCcM5MbclE9/kC2SUStjLar+1SdwH
iOpcq07XnFK8YX4uZ68ZCWCC75GNg3IFlV2udCU/Wlc4/KC7VVTRTniFaLUcM/u1
dSAHiNqz8WILumjQbd8HOYFHalVuyzVCOQLqeqdK3RInv3waWjN/jq7B1qPg+BjO
vuXeh8VafgIkO0+4/6OpHUEPB7ScK7aKSiCWdKqCU88HoRqeMkDu9Il/VgQrq7nq
ecIH5c1nkZ2sYmsDY/j1Dv/vhFEzi2AEDtgAqDO348fOj1jVWLRvx3jMrwu2HK68
VHqH5kinqquhLshY2qJqHLVh0ClNzLPgqBvATmQbsRcmPxxRXp3Kq+sCYOGHL8yY
b1522LDVJo3NYvRXV4iXo4sT7ymG7eJUVCvAsgCgdbUaApo0GiMObGAYUenyyCcG
1M1lTjzS0IDqDWYR0gcITW/xKHLNKwEjpYFjnwyNa7tX6s81ljoXAZw+XkfXdE/v
YQeE2v+JWwW0Qdl8ryMi0tMG5aaHyeIbSVLes1WaNA103HRkDX50xcwQ34CyE0QI
9YwyoBvw1fqakg8PbE981+KtRtuDBVe7P8CoL2YSiBwKj4gLMxgdUWb8QuqQcxxK
sskSKtZUQOwNyvA27oJGIRzlH180xTmk+83DNccMzSJ/c4QrXFEUrljOYGvYh8my
+0HZ4hyXqkNs1G1GKamtPc8rhI7wY/7xMLaF2dff8lVbavFeTO6BAFs00vOA2peU
EzC+D/bpDIGWbhhV5LCrkv4Z2HZKpbPoveppAnjwx8UgSPf+8CUKcJOua5eRFMzm
/w7oNGkEnl/BSqtS3rMxYQZdpRWb3DV9qKDJ7tMtrG/TIrKaNHki1tTVrDnmLTwx
levxjEts9QpfuPPFxlp3JJXxxLRJwnWGzyNgs4Vp44g6nc+LKwG6MHX3XRxg36dy
/H4eQLOOuF8Qp3snqkOZsYErFAaHvFouAWfU7mh2tHoWu1P2TEw+yMa3PG9LGyhk
OsWZ7/zLP4ms6GcZcLjMHT42BasWPphS4OnJqXCuzBNqcksl3iGN3OeWMHWcij9O
yLQQiHwUJZGHwenlqFZeIJpgLXv69X6NEeEl38DKmt+dGV/jY3e2uSp8O0EQDnv9
r2pPZdcK6bPSkGgdeFToS9zndGW9rPBhINLASqwZajfAdg81rj7Biim5ZzRghRhY
fBHzRHzMVqgGuw+RZQUkYnIhI9fUSE8bfRKmC64O4FBvl1Hw1ZnopD24LGeByTI4
zE2qm4ovUu446goHPjUkRtmPFT1IjblEnVAnBUH5M//5ZUCHBNBsI74CO/syWs5B
yl1vnMUOMrLk+SSlAHfEVHuMvwRawVoJf8wj6iNEkd2ZhjNpmCPEdlyFHKPYgjXQ
MJoIIHhXB8JfqIYk6QoSe0/DnsP6rvDjjN5/Kc+okPszLDmOY6H7/Ji8b/hVpJuv
GAe808Jx8ohuZzAZfZYrGfd4iOIS8D7oDGVEOBzAqOCb4PA490XmL/wVKZbgcrYw
92gZCJvVzKMBwQNRYwvdBOusUezves/nR96ueHQNtYJf12KmogJTmVZ1vF0hTPWe
Y3++pCETsf4fsg8VUJmgMDLGDlmbpzMFyT7kwTwQ2VlwARXmYoBAmTSS+WDd57cz
96F0sOpAPgEuzdncwiWBcSwXGaxj/Zgp8mBvPmCMd/k6god4Z5hzAQwENRXM8WlS
LooQEh2LYk94gE5vBRcKWMjJz136i94IiGwp+tTac81QimxGiHSiKfX38U95S/OB
A1iUVBL7JPWWlKXa8vR5p/0hMfAfh7JCImdOuc1pD4k1QtkIsEPVLlZpCvEhwfwB
LFl2b8kGPVm+Eqe94YHe9HyWwGlW7vtx26ytCQfe+mT/BsLDYDEUeuvGoZK+yPhe
dNbtonomzkZojZtM3D5o3PzWtRoyDwSZvVlCmggIgHLTr8rDQbmfrgR9Shohuf5Z
DXS33qIMjzPQCvQSD/8i4c2W318nf5mK3bZ5xiPfHkcchtI2WEgVJBBSFHttpjRK
5MakDoZ827x/ar/9ZhSgWeyXMuTl4SIrqQJuTsbbqujRU8X/0BcuNBlxr2Au26wB
o/V3OwomZVRCcJag9MyzVfqXpbpGWq9B//HlGLRpA6cLCFVFX0EAJLv/sv11c/ur
UG6QJMA2I4CBjJZtvirXqgurQdJ8h4wtBEaW5tqVdAnq4nrTKCa7f/zjqIh4ciay
NNlL4Jb94VnI1y89Se82Nmb2JX/psxaAcs6f4FUXF8LM77KP66lOGQP565FGcHXM
HpRppHNl68w/cMuqhSEgd2nhPp4rO1exkBWR8yNzfNwOv8aWWRUMnJjyy95Sho25
S5guA0jR5jQBKQQYEa9X8+GOCH4QgfRdi8GgPRvZycOF0S41ALaBKWsjaz8Onhs/
HyOOF9pG2kW2ndX+dtb83UncmeMiU6GK+FJBr+LDbU3ykjP69xr2TkUWYsQAtpDq
Yqg60fPwMxaSKfFy92FsuyV8PzgHT1vz8qfgPRxFLSTS7ESA/w05p2++sUMzJ/jC
KXb7xJZzv81zKYfDHj3p1uec1WMXKtmtWNiKUzqA32/Nf5QDi8ex8RFgnnZXSbU9
0JyXZbbNsF5YfMgNXI9m8Zjz5XTy58dKkgF/XcdVPJVdSi7XPne44JFwgwul0svc
rLu6XmxghWUJWuFV0TApU7EUi9fN/ww8FI9C3EFvjiZoj4AKBVNV5D0PXe+0KhMD
FmOA/jDgX63WV9J43r4qg+Gx9kC0rvZERp+GKZ5OHklgdoHKLDrygpdGvhGSvJw4
dnDoM0xRifBHPZ8/Vrqxky3rhNNiT7odCd334XATNlzwHskRJfV2Rt2TyrS7Aka4
Ub7bi+F2AAAMzejoGbKL2pcusWfO+uJ/YbIMBJVkwD8ZtvzEYAXy1DfwWN5WZjpC
zIl3+2KjtX+91z5pNVeAdy0u+H/bG2cW3dRFdsXpeNPlcqa3meplWkBICV921O5a
hy5G7xa2AKzdO3iMjTAd2JlcGKhV4hM3+dH3l7JqVYvwETrwoH8MRRFFt2niR6jb
WT9Vp9MJp866554z5ZpSwPaxtwzw2NvxTfWvNtWbe1GaxNbmE6/rkVdOiZiB98BT
oGya0iGszegF2m5Sk+4S5cYIAnjwvjBdsvvDLNxUB9XPaEYJPT2JFbsTDzclHxz3
bKifE52U+kV+Uc1da7C1wcOWn6wqItZ1+9N+qJpeOZEn/e+jxxrL59qGu+h11UxQ
5AVjXONY3F+wG2HoA7WH6HnA6K4GFJEZkwELFWorepYRYXhZUuMZIpuAtjgfjyIK
WxdNlvNRzsOAHUhz07za0wnB0hzpEMY564Cb8xgaxHtluJfIbHsHgfC87LmTO+wo
9fsokb7PLpMi6mkqZ14ifK3zVwSLv7OGosPWziFddmLAUI8vD8fUGpyIJrmPHWzI
1SYjL4yfTazRdWmTctbSiwm6C/AGxtfXVXH2z0d8LV+Na1zsStbhsyRrshOZyDwz
31M6FfpG4YoNX+AEr6H0D/m2iAjKQh4CkLqiIk9rjUE436uXecGDoaDuksECuNFl
itpUTv2WMw2SvXTbq2ma6Uw9CT6fu/P8bVvtBTvMDD4UGJSkfq0AarxxK3ITkMLY
WbIn2a3TZi9OYbXWCPxryOX/4zSe/mp7WgBTwhjnNiFBpONf+82kdke5gxGNZarG
bf86NsPXNAKv4Fp+9atcJ/+znxo4Qe6r0Oo8umHxXvahZDyDcbz+URA3r64rYMct
sonYmqtXsDkQhCWgkKL0ybLszGtaIoyXh37YpJT4Idzu0InZMmDhyCMpZ0Tc/E0N
M5yfKOf1Tp+QrQZp5CMsRtDJcHWPbtiyhYoQK1QuF8GFA1CIxWxDjRyFQAOgZhxB
bTyZHttITocZi/lOZ6qmhnLLyS1eYp+wciHEqyjplH8XcNgWniU6n6bWcl5aD8yq
/cZqdQLuVLWJchn6xiVPpqjeSy53pkQmsHYDcWSRXRPzlIBVVxjw1y7zXPo+060+
N7u0cLzVKS9EnypPqVCWz2n+7iw2pM0XtIeY9KoOeZsw5NC+Mqyq3ajn+BKXBQE4
qVtStYOpswcf39G4FwslBMcTnE7T3l5fdRutnYsfasg/Ab1s4xS2K3a0tqbEejoj
dEfg/8WuyyE7DBP7kwEK+fk1XdL0Hcn1uN7rOoHYDXu0Uvik8QrxO6qUALrGA0/E
x0oymK+oTFmdzkawgUGqIKLQ0fXpoVRA8o2/kuLnxiNs6nYwwM3l18DnawrCYHXW
dt3ak3B5Y3Juv/1DiDzSkJLHMcLtc7qfan/OFDR6ZIyTY8KcaSw2Eu2Us+MvH+yX
vFE7egVsQ4XNLuxBr8j+5V1rroW3i5TZVn6P4gZS9d98BH4H3/w67H/oP6g4xKCY
BHTrp8h5/37EoYxIm+Mbje2yni5E+zXItBIFahQBmCAnCBr1vZIkpgOahwIMK/fL
nC9W1QH8PoUnigM95B/qVnR32Ej32Uv2irueKNy25KbzQj5drS6Xo0jDNjR/E/54
WqlS2AQ6rFJEBSZmiIzgUQGzkVaYXkfXSCkkzMr2rUwsyiXu8uJSddalfxnLD661
1jMY5no+nbv4NpDQu51L6G47jthXgZNf1WnSxUy0IYkIlKl0PmswmgPqRRIYbmoW
njp6ba8gDfcldGlVOqYpcmwS4TNce6tBiwNNLgUqbai2azX+DHP2D+Mp3t/CK7IN
0cT0KPre1i0c1PGfZboOMQ7IF+BMTJ1NR3Ykp2wblZdoDXVenHZTQ6NuHYxpS1zt
pXEhm/h0RYLJD56l1zSQymqpOGVCQA2OBmLn01GcSYTpGrJkjKB+naR3u3INfGjA
JsG/IOt8/fUawxedY+ymA7YCQMXncOMumgogPpeIBsm5wOW+REhS61dIxieGXSGi
gOaHWVR0oVlqYW+YFxOWEaCtY7Tw7dqf5/WvvcR2IumvBspRIoUfEXdIbT59xJr7
AongXHHwOSMuexIzpHnI0rZ3gar0pbihsb4EiqXPIcYkGf3gBepib2m+VUvA6W+7
B+3zDTszJkidcei769U6j9bLe1B7oBB+8w8MOyh3GUuW0Why7Lup3niuG7e6Xxwq
oc7dg9x4gzysjTpfU9pnAjXEVbv9E/Krp9uvU1zEDt6nSYl9+T8TgzO3xa37/z7F
0NmMST9FZZ0zdxH/Zb5vVWE+C71EmQFT8jtQbWEATSyqIz0nPl/L03WC+YSr6gyR
lcqUDGN0OXKUycfKn4o9ay2xLkt77K806bpUjvWjawNGZofl9M5y6QqJINDM/OWh
R0Qe9akyBXSldH+i21498PsmKXOu5WhZ5iNVMhGQIKO13lCCcTHABoPFBuc1w9Kb
smG/YfH7gTHz6DAct0PimmWmxqbwQDD88MgdkrzoYWq+2gA/8zJF3IID6N3e3NlM
1vOy1cV3UJvkIXxhW8RgVr8PP2wwpAIBusY5Z5dNdH8pCOX88VzKC7kE2d/ipbHT
KdjEZWqM69GSuf96b0VW8Mg5WkuaLpuWZq+d3o3e2CwuqLtDa3bqJoY49fx40iwR
WqzEawG9AlfrhngKMpEF0If7j/Qs2k13uBehj4wT2pwz3hKzsw4+8IkxW/6hfEiA
g1MvxiKFQbsu7L8OUPtOR60w2puOb+d17j9iPeIRTrj5R/A9sDvaL+tvEDKRFs5s
SMw2sg8e5C0NZXAb2us6aZKC1ywtzfem4p4ih+AnNy6QcuTolB+2FWuxVKKUAGp0
y9+xqp4kf/exr9CVrI4bWuj5Ntj9YU6N7RPq4yqxO2BT8mxRhCCGSU3fopXiLI2L
PM9zEGtzJwBAxbTb3gdYkhoqfzy0ST6pCkG9arNqhrVuIh40wUb1CnoTj4XNA9O+
p4AL1ZVM+UKBqFubEcYbm37yzzJvHZOC99eXIp+GfCLnPVd/Qz2LwSctIy56y93f
XiMzpq9MasmeYHNAeB4ZrwLVWhg1TLjQv9+H6c55uIU4/3X9UQNH4gghXYqbxLnh
gH7sxEro2+Cxyv9Fe9sSYuNuLjY37YclzbPKQdU+m6d1vEB6RvxO7omObg/iN5g+
glA1GKMxUTr8KFnMnSAnqSlrv0m2mrhr2Z4fRvBzlrMwvJfIeioURF0kTlOD++p5
b1j1zrMSnjwJ4ar5cYQrvEgbXhOjMwy092eJgiv1h0Z1dNaErR+V/kg1GYU/8TAM
LzHaWwRIPNuMJE1pCnEG1QH4aQXjE1sUmoCkKWUU+d7Sa4g/9Y1RoKHHRAyz4xxo
70/w24ncKOyaL0tT7zQS2YKzNaTJKmSsQLXGemqIVRf9wug1Wo1PETVsLhWpwA5B
3zhMjstiRIXoT8RF0XY3h+mjDPR/D8QT2oOR28W4pCmDdIQ8q3p/Kzz6+a4fupQQ
f/FvJhtjv8NHkQcWnOdC1SKRqHlFgE5w6R+0pfXLLSIrPPnpxmOdsztdkiH0Mu6+
8e42FAXj9okiuvf80F3BascVoWaVOT3s9UGodZoc8omb9DA+uGmxlmqpQDmzYKGM
uGy7RvlH0EVGeet5vkW1HCtNbdi07dHTWMCNCCuwemlfjuFd5HmD8oPpuuvDGavq
ejvQKv2NitrhdEWJIuO6hTRER3+ElrRmKr/B4bA4aI0qKllpBlGJ6it223Wnfc6x
XPB1p2VvfgTsK5JXW3Xkv9wy+WZ1KGcl78JCTaUTXPAYzzlzFWz2P4SNQMHKZCSi
wn+TEY6LgRbuWlHvhXcdB5Ua7XuMQLw40cQZpNNKB3JKxeuEtULC7kzr6AmllhSE
CbQ2Ku8uk1/I1J16StHYJBL40LYRlKAqTg1ojqkM4ceaHg2+OPLOE+5thFkVPVgw
n/QwDYgs3UJL55QWy2U/NZwOY0l1AwtIY35ABmsNpCLUbX9JhB8z5SBjQ0OQCfOY
JR81R+cHLvgTmt++YGa/A/53Xi3j4A2iztJ0BPY/4YWofcCPX5oN2lDAk/Th9tCp
zXiDKO4wyQlLCPAS2dZxsJbS4o5ovoEKXAIy3zsgtoYwPnRKY+U3xSOukHYotz1v
TGR3bkhZGL2Mk5a+jBQDZkIkpsKzxMpKBBlSFXhQClVM+dIh6egOQurFVwsXBrnM
3Sx8VjQOyS62oyfoL5wFS5rVOaBaGnFGQDgggg2NCMw/XH+/zF5230VTAWE88p3e
f7rYS5I7Lq63IpMRXA9V9khzhkpAQE/3czZy4YcFoSqvdv34hT0SsgWuKmZLhli7
RqSKGS/zl2RfvsWCobfCzdim1lPsbEeo2fTGTBbLFcUxqMgl4PSJMKoRLdDffa9e
VF91xiveGS+PiI8fp4wr4rD19JZIUAVC8FcK6BKPfyoyp6OdNAz5NBvejkEosPio
frjuz1AsEK0TCOrAMU0uRRDinFgEVB8HEbnhDHJ0xJqEPzsX730r3lbxifIU97px
QjQEBVr9QsNvb/nVoK4dzpLIm4emXzVrneVziiZK32SBIIBFWYjqpbYecK0aqUA8
bSjaLwArtRMpMus8YieLaLLeiAjhMSUTpb+/N0JnoxRiNqeKSbl/Ai05abacoAlq
oNaa5TDlKYss9d8hB656gDC6DvJ+xqCc0TnhhMUX/7o68Uus9IubeeX6p3yP9VZk
coKHqdRK7ysRYvbztBU8L6PM4PmBRR6v/+Rq+drdK8zohCgzBZujMUD1Y65s6M78
K9n5M4OOV2sYSQRKzmMUiOzlXz4S4JnFyiYJmz9nmx0Cxq1sg5/k30WjQT+ESMrB
PFuRBUGkFmx/5QWMn80BzZMwYUAbXETA0P0hGw356L5DH09gfKjOSV/xeEmuvsjO
trO6Y1bKiF+qpageXIpQ7MyaPB8u/FCKujRsn/Y5+oxiZG9r59vXsqOCBpHHCDqu
fqb/9kB/eCsPrMTMxvPAD6GbDUYtQEHP1kU0mm7Xu8YfNA/6Fc+M2+enOvoxm3Nf
wGl5mPtu6VvtFRisomlwkVaDi38KY21qy3JNmmAO4GQZ8VMwpF0IqLput0O8+Gz6
hFhuJhLuUe5q94etjW5LpzRcnXtboSwcAdVkk950fT7iRQKs79wojEUMG1pRTkGb
EgkOdLjmIuG0ZDIyix7fePlffDiYwJMpo+dwldwx88EKbQeKQNqSOWXifkC4D28l
BE5ryEqNrBNxbZzFAaTH9bgZC7Ancv+wn9w5K+QHuhWkAWP7Leu0p1INnZMEhzcR
RTAf6+Gzt8E6BrXvxt/pmduEYzHeX2v2vNd8KzfLvxjBQzHxV2qMBHVsLMpWLRbW
Tx4jFOWfb22gHCyLUtun9TNvXMMyPLUpncqWiUSuvQy9MIZ22kj1SgE+G/dNAt5V
mZdT1I21U2XKFE34yKDkbs4mU0At+OoqyrbllKGB4GVsv/aa7Wh38xfzuvC/0uSb
+ZuIp3ZNa16rfOcrjq2wLyt8RRKwhNuOEnEc85LvWiaOwNGYA+9mnB3FzwHNc28t
Xgtiq3BXpc6qr+i+qP3MTrmjWbEbi+eW6x0WRvhzfbG8aajKLfh+Ba5PHcNhiKbn
AMT4eO8Ko+DSDi4wb5Wn8lKZHgxH+BI9gM+CCIM+9qVDReWLSFFshASOrrqEw4QO
LJyTmLDYprJQrykTICT0MtmC+QHzUcS+X3We8Ag/XcpomHMXlmowKWNgUMN2eA4W
K+UfPEKKP/yda8D+RnEJWfrSd3MPxwPFLCAKsccvum0HGyou5eCTq6TlcTuRdlDJ
yiqhWhT7jkbH3lfFMe1LBYFs1zm7POai+9A9pkkV+5GSYqubGgPifFMNgO334YDy
6GAbDl+l/fq3U/5W5+JOgIgidRSrAOMdaMzxmuG4XLDcvnADM52pogNeRMhB9nge
ZfsU0Ph7T2J0dqpvYre/DrVVGirJxRTJeglalcEGibJbSzSOqc0xHkvhnuXuOAEl
2jd5oS3epIe4KYJ9s0S2zLwdPQIEm6hNyeNuA+0+sOWXA/lMulyisq26W5eQw19v
t1HZZ/Noi4LvgQUxA/befKH+nx9AavyZ3SBzeybsLLpPJGbSUu3B7V+0PaMXwhj+
ZethTZ9xKpZwEbvfS7xlAerNQ58I4Y4aydjEPD0M3LJZY6uH16E/WAh5sr4yXepW
6SGVpptbztwrlXOBO4mP7dx3WSmxyclu+JZeo1ibAGwfu4jkGEorS0sW0lS15kzY
X+j4PC/Wj+qlaB+TmsVZHzGODzzTvWO/qBRNQiX3hKW5VmUCsuNdgwjbucjvrQoS
Imk3WgoQEJph+L5OKz2jtj8a8emqQK+tI3/UMk79SO+aVeHzFUQX0Hn3Uv6N87Iv
c373hNSwToj16CCs4aESZbJWUeUa2VPyLq5oJis8O/8B62DFDhHlEsz95f5i6m4i
Azk2WYlFvilh06oM2s30cOLlAoDr15sUmGjdCdvmDlomYxHfiHdLd5M3FLt/Ftnz
Z+ftC+kaBN6477ZgRqclgFjarUwd0wKOTaUPi23LwPbjkEb4zB3J/aR32lvgkP2A
B3kfObTrxUP6pKP0ZE2BkCOouinZRfbpsrZd9+Aai0LsvJdUZQKlbUS4ND2ZVQ3B
MyEDjyXa8KJYK1+1IaYHcApUWNeTAKA5QT7KNOvDDsB78j9dxFJaoq+Yjh9b20nC
cx3lrSHMWVbYgceLzsUfO9PdAgtTyBrsxHz26XpLQA8ptUxo+PEnIcwIqFCIoU12
0elE8N46HuiBOh1P8yVMVRCobzQ+n7mpNExC/R6QnrG71tBjFKr85uCOFBFmWit+
bSlKqLpOw/avLnQizegxzk25teUy5+DhtRBsmCQRWK8hEe6SjD99i9vp6YgQuLTN
dHKTdtnM23jUYgl/AAmURQAkXRoxdmueWxJMKqwx0wJTSvZ9MmZVs5LCIbbVGrnt
rfn7zAL0fUZcMi9Wnt5lTRfdokbyVQuzSMOilxILMUWd3CeUMeBBxnTsU54gye84
JFMpTgee72WYJgZQ/QKZqSU8tN3DnpJ/ojxxH9ASZGgL6c2U0CA42J5Ua1RN7gdA
js//JZzLAezJLrQVla0iT/vDENKS5ft+IuFdPKpGgJBeBz6516ZcqnJrj5SwsWfS
vAy46Ezr5olPTO3VZ6i0q0nga+RY3pTdTkuGOqJnbUx39bu2Y0HRFXybzKqsPKa0
mcRUUPQpYZAVDJ6gGwNsCWzGBlnLPzEvFphd/Jcs81LlnKyIs73ERqk+icrTstSR
L7eBp3r0IbDZg4r7hLkgSnf+tM9ZnxPyLey1U/x5x2e4Ea/thAuUUe7HQeeu3ff8
W+O1TGuACPq22UT0sR1oHWwG4ebrtCYMiJh9kkxrxsPRn+dZqJM0GzT+E9hrgmRG
C0ImvkRKDOL9WXGJTCHwJJBKkULjyIgSSB8QnNitF6BkzQyrtx2sovRsl7npu3v9
gMVDHrssTiL0losVZq9fdXcADCP4HDwUO7J6WljSPo011TXMX6bbOahXVXq1Kmea
T/LzREm9S4fTzeGLvCp2md8tkARDFD2Cn+k0y35kZX20uNtkOaGwaXPEndHvUdvd
izRgWZU6CLr1jvv+SjoRDtMYxL7YTkZJV3+mB/JbtZ+KvZoLFxKrlxZ0eE5ytM+F
sMGiXP9Y2i+WwthW+puASShzioCGu4+1vgU6CXjKIkAC1GfT0WIwZkHFVUrsHDsr
wRcTC7bCRtmBtskOiHC3U7lMo9rmq7GTa/ULkwELffsX6ZnzsKpfnTLVHFN0Z5H4
LNFh9KVNLpw0yjg7P11+O11YW45So+u2VLZbvg9lB+rDtiY8mDmjbZbZbtp7j51l
0svGjezaPIsFbiz36fvWorD/np1ipqUal7+WJvWlJyvCFTmVbgJxoEhf/mtGZ1V4
08ctf60cXOLSMqjahT+/vy04UnjTXFyZwblEesXNnrQ/Jnac6dR6zi5puJrrAhuB
j2TY4tep9dg78+4tjxfHsMLVGxo87W3gShTteTlcrVYp05XF+kdIRJd9/5/Bdg0C
dnVVlVS5k/QSJb7Vf8DRum6AotA3nWjDd4/z4RVLfh0rEmjhl4tVxaYkY8Ft0CBC
yEP14yhiq/EUpp7azixvOX1TcxmYH0ArLCb6ELKVMEMj1HE6fU4oToBYpaexJHhw
+UeigX6lhDDBQOutNT0hb3VQmdYgcMGxMj6VltPwAOzGdk3E4FkA9vtWd5e57kZE
OKSTtnS5QN/5UFegqFW34JxxhmfMHlP/XZn4nnL+ptfi1wPGDzK5/+b9bxv1fEY9
0A0zAYJEBsHeeDMY2a5HyYkGlXXTI8of5kLL9xrMhzLSHJfEWz1ppCXt9Qjm5CIh
h6Katuz8CroKHzKO17YJwYCPDwQIJtRihLOa7FP9aNZP03CRqwb/LoKVkxINSFlG
iMiI+rg0i3OTDOLn2HGYiZZwlmGwU0s0oC8DdzWV2B1zOX5IAx7BqJK/he22JlW1
GawBxu8Md3hEiGw+PDRztEBBDnibYPpAqrZ0nec8qyt8X0vDSqAWrA3LWc4aSZGa
hrIYocYMP1UZKHimKK5JSU0gt4fQ0exanLPR7ExBkSpzW3A5/fgoQd8gVcQqqImB
G6LSHXx+zuTnkdbUmaQCg+pBB/N93oYJjsUWCMb/Uk+VvSELmXwf/aI748lIDShz
ENFFOOrUczCTwgwClLKlpwxkjBK/FseidCaF0584ESWk4ez7A7Eft4K++cjvUql2
Cmtwh9VDXb355BYBJCcnLhK4IRkB9dA1VGKxmuKeur3zg1mLFSgk/VzqR2NHMSTw
qMtov2lQFxWCAWKSS+ebcRAoq+aKTUH1R3ieSm9I4X5ph8pADRNy0rYDmbeDt4Uw
Qrhcc/0XnKFknMTErIrktBKGCTehvohQN5aVjASdjN9IDr3vkUqKE/lTV7EnTDr2
sE099t/1kMev7p4LcveiaZFhxR2X1iupqVuZSt1XWBn24Wxtaf1tNm0tNxKqnLUc
ljXPrYKHCrOQ3gapQHfWosLeQcojQLPcD4vl1MHcM2G+vZ9JBXz69aS9PoX1KY14
8pmxipZ0+8byEW+ZP+jPZDzr+eEDcshycMvHYQJ4ao3mPAcyO+3b0TPmy3ENQ90Z
WwGqwgfyQafbfAHXifhLi+l3MKTnqa92q3kphzigGs6Nr5Wwlnh/xEWy4qo8mhcX
rDXeQb4lzdzaJmdmG9sDVlZwnr/0taHQkk7hxQeMjN7DYnzY4ijjCT7XFqvNEQF5
APn3mpgcSb7Rii+aq0NGdLo15G8QLYnfISfWjJXkc4Op1BRd8GW1/3jSNq5wVzsq
u42/TRg6bw32HgEeUroRIq+d1lnN3ZOBNu63dVuTJzEvBEFIojJwd0QGF3GDdvoJ
Gm5FLs4HfRs1qPyu9aCaeTM5OO2mH50bJkZyLvuMzhWPZQqqJpeywYHsXJLwqBbK
lzbWaGFvUjRCAv13vMox3+q0WHDFORGvC/RhVzmShwh2kexf2Rpq0iF3Jp6n27hG
QWMSnGDSAM0Z+wPU0BAndVSA2YcQDJ+LM20Er4XWVLEk0t+fNxLrfIL5un02WJ6d
nFSDpX3XVpt5xiCMPPI/M3ILrQYM8jtp8z/ev4a/5s+QWpv161i5bpPVNKW/Cp4M
mFjvWNMEnZXqfxgr9A9syuhRprPHdjNz0EYYbnrF7RI8J61U/svWwW2YF3segyAa
2ODDlzc30J2ztSPXOomrs/Yo5rT4ekJ2M8CCQfKcS/3avzPD+I8QTuhVz6quHTaO
gEVdKsZjj9GjVb8etyEdUO15jg0Gz8EL1FLGgTCj9Er5hVDVh2F3CAJ9O9JZuZht
G6pUa5eUDqRnHeSyEYij5ZUD99YCdWz559HF24rkm7+EnoxMf/lNxAzTyIoqTv6y
Yavyx7C5aLsffP+v1p5G/iDfiuyd9YheBjJJcBjv5MqIsoV3lg6zq1WI+eH3bB3/
6eGF3eSgzc+LOPgRtX6fk4aGfnROLw/ZymqH8AMjG4xyqcG9t6//HjFQfwOjjOLH
mBWbnXHmtP3ylZxzm09BqYcLyEzHhxCJO+rQbXa+JeXDbOTHJwBjQBkH4T6URpx3
b+6HB7AoLpd8vz9jX1j7V5tTJtumg6wu0N/o6FHw/vY2wl+S3ziUFfRJDpbSgsAt
L5bBQG22RHx7KGZCDbFPkTWAeK7svCn2P2MCsmt8XTNKwC6CkCICxg574dvji84t
W7nMJKj5zTRj5HGvmNwhF5xFouBZo8TYSr5B9DOXj8BTGVTq/vai+TA1ZBZwBwgp
WpRGgeHBBzbPHYQSftaC8957DgZjfMZxYjvnHz3UALgmuERjT9KbNVBENwqs4j8m
z1m7E2lAyPfbdATT+zadgw+K/l4ew+GZV0m8cBJC2Gx64nBPgWAD1C+2DXYH2z5x
cGv0V6RYY+/OoEA/33DwbPaUVo4fNzHTW9pQu738wPA7iAWZ5YclTNxw29ZIZoRQ
kAled1xJz0JttpJr7xSSW4dYzpeJz9JRIs3FA1gwegO8CCX8XYZeUJHLkbrNzgmt
n7WbYpCC+5g8S0Pib1P5loFU5s978PNzDVV11SaS4+/ub3kqe9jLqJ06NWZMReqo
ROQ6goEowlIaP6QZ4jzUkhp2Z3kObAy1NVSDNBZfZaqK6xjlLPJrVn0ySy4hhVan
AfC0qr0afzxX5bXriIb14j2KzAgFbdmt7r9Up+JzdiMiWA7I2QhPBAatkKe7+NAE
9p4urVWqzRTS06ECnNIGo0pRRws05b6pvsi048p0kSWKtlOQCEoDNcLQtq5DNjas
uAaZdgMx3tgQtEZepUesxgo8MhueXIicWHWPoAEcq0ZT4dYKGfOBk8wc6uPLVloc
L0jTwl6U/rs6RvARavZWsOwl29wF4567kdP2UPyzi6DDVGc6s0xqWpHQMiwssg9o
3HCtJ0OKqx9t9cmOOBN/pk1lOi013w0sUzHZmtZFJ6e6ht81mMFhR+NYMvyR5oNw
jc9BoO0P4nZhZ9Plt5h1UKS4sWADUtfzL+XFfbeNnUSPGH18vaN8fgdN089LGHO4
PJ8lCZLvKWVHmjmfVuq0BxjWiJPxvckarv01uOGSgp1z3a9LP/hfxoXVS48sBcyR
jZ4QljVryO701fbJT5aKf+zDwKRxRldTa40TGVFU1JzfZMDnMjG+R+hgGIjylXnm
659eR4Eo+QC7jYJovmEZPOniIbUUYQq4Z05vkajVtmRL7QNsCpszqSSNY8x9vu76
8gR1gw0QIL05v4weG+MCYXY0/0emMOLx82ZOp98VZ1sBYPazjhyacr5jNWkVxfGM
OBJz845KbRkfAOni7P6U7rzbq9luzmgTPIrubJU5l+TZAh8hJzF+0sLgEZjvQcV+
Iej3Sc8p4hm+di5noftcK/4xGp5euvYBGN2jcKkRXbYIeWB2dOu2D5vqGWO8zfDe
pBSp3QuTvHdJDkVewBkjcT/rl+hxnBV8rcQAmcdOzin+ePpbXBBtEukVqYq9aQA3
vUL3RqbFVX5s0rJ64bfSy/LRLeG9u4Vyf8JbE/yq6H6qFnJmh5/qIK8TdPT1Z5Ki
i2GMCwRtTnddLEP6aUpLQkbdwkvcyaHbcSUFU2U1mbUH+wKkE/vM9U26qsZ3HhdP
k0ZGjel6/1oSxM4iAP7e9Xt5OVaqUVZiHpAiatoI4L+qRolCDgzByr8XAospfowX
Y5f2W0J9haUNY51komjOPohAru97Tojb9OE7KcxHILitwjubU3jVjfnjVqxxXqHH
cu6sFlh4+VRkOGI+vjgE02uJe/Oui7KkCasjSLimTrAB7CZZazqZWp6U/AWZZyM2
JBFLQKUiaQo1f1gz60fozXHHNBZJHHlOEWGYF0DC2yCjrUV+wIA8zV6RYH37onwi
/3lMA/x6MJTSfm6NWTvhkWkl2fbfMJFNl//c5c9E7H7vBDtsazxEGiIfOZXz99ZW
Ava/pWSw5YHaghJ+o4pdO9un0Lfgq7puCxC/scf5r2Nvk5i8WZBEzUJIDVEqFuxv
PnjSF/hA/4GfwXCp8/w139Ax4HXNoRLarTdsG3carFbMpD+5I86YgZl0MF9f2AXX
R+WYSiyMjtjfN9wxlzQHqXLYM+INhuLuFhgCkmrbDYbeBXPAJKI/X/FeKfVNLmbY
8cCUOKHJdNsRxYARO29xefK1609xNKoYNuzW3V5cay9sMy2Aggnzc3r1UwWJjZ8L
2OC4pFAHdFkXLmx7sAZ4PVHhZkBUqPhO+bXluxbQuQBCQGtofDLw2bVzxNDaFIHV
O6VYtpHazYkgOE+Bz0oSaWzJWRVG+sYlK8LrBp9TnO/zrxyxlGNERdGuESThCSgW
TynzuPWw/Pkk1t4t0Faw8oegyz1WktUqFzBNLD1X6sAC2qYM5NsVh8NA8QXw+W6K
48PVl/0KZXTHhf86pWPXIa2/7+t6RsCt6xmvkSW4MaRMhUF1wNadcojJwVfdagm2
C0n5Wsgli9pbCDh3m8rH9WOFXwgVz6j70ZvhJFlvH+JX+WmWS1rvvyTxwSpQKaUL
+yySMmi9i/FmZJHXBbvNGLZUBtRNcX6v0KXV/WcLlVkCCvQszVMPEdzb0+Ir0tmU
3H1T4hslOkRJXpb/pZV1Y+lnnTeWjvaQYHcn0Ar2y2vcwSOwDof7XUTYtSj6GWWP
NQ5Pw5QC1iBFR0ZpYhoMn3GuJBgh1i1VgPVJDsC6PYj0Me8SIq2t3/xGEYHQmK6J
+3iS63ABxgnRPHO8TgAS9xFm05N9FhS0mcVoQ35Ed72Lfuuj1B/3wH5hq43H/0Xy
QOAK89IQ5lvW8LlEaks+gAzDBkE7TVn3Kx9lJulKcIv+ETiW+jotuJUSFKTPg6Lz
aZTQsAm943Z99qBfndIhq9D39o/a+lf219m52/s0BYcV/4FqPfie1eMqo5m06dlF
2vyBYv9WPehsQ83VB3N/FzKjjZZDkLo+IKJSZnBBq7zwuDod7SB7AuzMXiaEjsVT
SGB+D+vt7zJeFayO8+VUdxeo7RLLd8h8Cc6KXrzlTe+sOdCA475zA6MRfBNfzmqa
StnbxQW/cFiq5IVyFMzKf3GDDmymszYVN1pJoRIZA0hwdATC3cicDsyGnjIeXAVg
BzJnK52h58zuMuPva49akL88l8yJJQ6mXx6NuvtvxUskkYcxYdgFm5+Bmx3cTFoq
o0mmMa627wvrtt4bOG4AGF0qHkrXQNAiRMHtDY+J8z0WYs9nWQlsoAy6hFRIvwzg
pDNMRjs6JOTW3rglIMcToBSOqG4W6mzXCKx5fW8DjBaruDzOxBZbOQEJwj4UDwY3
Jb4C+wTbaTx0ciLW7CVCfbQmHYNvRUFBPLd4vJAXPHNqxILxoft97gSzdCr7MT5G
oWoq26psB6PHnkqywytIkjfzCXM2JBeuDSaDPehOrCmzaoE5c8ypIBuhJxW4Eu8m
JFr4oo4GTyH7gddsYjkdIPBM/CX+U5s5vuF9W5JwUbK/7feQU+WtBeCrjjsq5+AE
b4sc+5XvA56UEgVyolfRkdugjV7LExAE38exlA7jcAGCY9p7FvcIqHj/1OSS8XxR
BoU9HmMwdVjUo4QruqBKHOCFH0W3/92PluFWDE0wo5jr2zm0jRWcdbkYALq+hodO
0Z52fOBtTwtJsbJKnyL7jyUL+l2PEwBHHsYd9ANgW89r5r2z6r156eEvnAZKfEGI
Zwa7smHYKyRHBfDywvaSLRz6BGn+yDr0va65QsTYv072/cTBYGZEPDImbt41/Jvj
u1D963r4FZKamHgSV97EHIu9aU4f6nnXarI4RAGBfkseVocDwnR1Ac4UUsjPoOy7
L+tji4VE+/w3+0ttPGQE4YQZF2SrkbNm5MTV2gNiU2EDshUQ4hNVFG1ybCq0sQtX
dMlSKg719rs4brRZ2DlTQAhjEqcZVeoOyvCoLZDS25j1x8uv2XiwpGsPMSTqz01i
wEcNaT0FSdZ+8lx8vNqy90ZkmPJL5orxdaAfdP6WMXkf3UEUUIvi/VjLJuNwQ8HL
maLLX34ZeQqAj01Q+YAr9ibExuh84zrGw2f0nzSonTBdJcmABFVwfMDpXwlLDNB4
2Rq0B7VLj2XSiNF3rByBkxHTEOFmo0KSdmD69aa8WulWlTALVWKIuC6CQOKwxTIY
VrtrJl60vZm1pDXKg/1ELOO/gkojNBxn/b8EIJ3Qw7YaAFH2K6KPpEryqwLWi2Ld
SkkWFd9yNo2X0bRd4wtLvrwrt5Tq8c93T4XJewCXwUW37AE+PLiLABrG9bcZzDc+
h4CfBus2cIYWqIkgLQJHetfnsN7VGVQlqmqOiSn4ZSVYy9fycyoprXXrsn/8+2i7
8/qBECufXROqbVq1tSiqPEakHk0SWTRxfevTKJTZDXRdMsjdXQOq7LsRgH0tp9Uc
H3rLhZqGOIi0XYl600hWlLdQUMgetiLWmaOofEXZfoyzNf+T8sYqzTXJGuMhObUw
4koTlEl3uTFLgp5En+w285R7HktybLVWOOwYO75/6ZNsHBmhTLPEnbJ1SVk5igWO
Hf2J6q5f7KICJB5LEaKtLeonqClHobRpIeRemIlyMNHGrl4Yq6x3bFhHxfr6PX19
8jmNBohJxJWbG1XuxBSamoaNWlM2fAK9I9UAWbn7EBtr15FqcqCuLynEjHvh9FY4
K2mhMItd/TAvBPFdgX0hgipafA9/YLwPKnZTgQctPgqlQngEmvdF1D3o2CrlwG+z
MvtNucFq+k73KBPM8nmZt8sbUkTqqaeZIKz/xT3TD2y1CDkQa8ayXqlv8w0VJhun
/jsDY71ZTgaS7ZhVDUFx662C7e6cpGN+vxSTzM9DVdMjmXtX6GNjVNhfKcAnmxSa
1Pe/mRlMchvnlAqpqGCz5HPX0hFSgLveDh2CpbuBkYJglMnvfWNqxWzat29/POog
2FDdiGF5vbxXowtduFdvGXj+ajWBSvQG2ZvHBz9IxFUHOa5wWu9RMYSYiVuv3wIh
JET1V+YcBUbngj0OSz7UgjyaBzcysdJfUP7R8l2GtOElPP2egF/SMMBQR8Lmll2L
/aEKpeLFOFwAX6V12IcY5B83UzXgB/DeCD4Gn/qBPKFDhFWL5ufnIRgOUHYCX9QL
CBUtFLH5+0DuerZoe0ps9NhQion26sxXHZZTranITebOCLaATLxrPtKR75A6bSRA
5jPtaf1gFgpgJzLAesWffan1xAmb/0xTlU1lcdMXMwd7Z/db8ZPaXx18407hTN0v
KjUcpaB8n6SuXmS6WBHn0z/SWpK8/QZHpZP5dFeaCfgEmUuVPa/erMSkF/3wApM4
EPjvzIOJerk61Gf2F9ooRB0dBq5Xz8lGq1zATWo85naRZklu9QJwWum0EA2iHg4b
YQ/6Dq69EiwcojZcmbt/qzJgW7jVaYfgef45s4Inz8K7rx1fTNQbWOIL3h7/1YRp
aUPMn4KmwiFX+WaBtDL0dwv1jrsA0YM7Q4nA85sSXI+7TRyq4LICIYOcRaU+0z8I
Rx+mRnUivIQ5VTHBws41nJW964hFRptHZZcovwBVqdGV7XP8Y24VbCcsjbCy2DsC
HwQwPtN5V9DfZigPp9SQTTIAlilSqJd7MYhoUGV2iYqkIw555r6W3ccoD8jPhty4
agjJ8gH2FKa1NfDeAGGStfznJQ6Mp2Xzc5LyGnhT2F0GRVzpmMfwwBtXagyYu5VP
JPsYf5kwhnNtkpxXGjHa8el/B9B4W7nSzlvysTGDLJJ9PxpLQAAFaZTbaIMNRVvk
yKgCohyRNFOv1xB+EawrjkRrlByJWYbkHXJGgR7aW3a5UxNjBSjJNhhIpAJVngno
oa1GUYnR73zr7SwawMEhbF5ydZKCR/0gCCyyWVTs05DPC7oG+DWHgOPmfpJk7RxA
XWys3YbP3nrdzt+eaTbCZkpWlc9ETZX+aLT+u3rBhHHY0jpbBnnSk6yBEJOUaQA0
PcQU06uJi27z/DErKDD1U471cYbRkYjVO+8UK6e2cN9i8ZFp3Ly8q3UEVMkhPLz3
u5bdQNCfwzDu0g5tAseEbRU+wg3YGqOrFNo2xjwjgDgw7L0GF6P+++cDva5Ag7P/
BNpfSjyqlH1FLtIZe11vebekjmfd4mkjBKbiQoZr0o3GoD6AEyboylM6BXbaKF41
fxvBKT+NB0TYV6J5Co025nIdgSS7Eof8ZWIwu54I/ztMDzdK4tmH+9UGc6spCuz5
ija4e6cDxyrj7I8OMetDoyzrSLklHAMcK5u7W9lIkSgyPhbId9LPSY60T1TpaQJ7
ZEjgE/xF6lsUQYPkmg3ksJyr3ZNW4Lk9ge1tX5rMXRis4mH9VMTyk9f6jvWb/FF2
CG852ndBASvpuAyW9Xy1v80q+CFltB0KzcgD6RKsDrLjuizh3a+iw7unTFO51lNp
rzbBt+W+Xpobvc144dwW2hX8MNAM4FrmOktD28/rfZxgF9oZO7AzRAYamiOnE/wT
gNYjEmTLt784Enu8fsbKBdiiHx1njjaV+WXerFyLe3lvpISG63wuh93Ads0DpRMI
1Or2gDwYmWhtAkkUsxJ3Td0RjVzFdEHbL/hLulSCwRonARsjjlx0fF4aRrjW7gFS
FHl1lZgD6vcROR+/UnDCepM5wZy43DBHTi3aEhFBH1Q=
`protect end_protected