`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 6048 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
V11MTbmTEZNSo/1VkQJYbSDi7CI68OHKf1JBrArXicPtuRwqz5MBDGg9QvL5Zr00
7C+r8FYhBZymEkp29lghiQB2heqIdtctB8DpviwcKkmsrgbtiMN0lXvbRJRyieJv
vpqFOvsIvcBcya06arlrhPgaiaBEUIynb68TScXd/q+M3OQyr+QX8W5qcD1lmoGK
FTf4W8t00vIyN/X7TVl3U85j+yMmmPkoPhTmPnReR+KTYpWnLbhHoMeyfQOgXFL4
uhO/i6JGIhPzjz+kbJuFIN+9Gnknw8bk62PvUngDg//BS7befjDsFaqknp5avVxy
WQ0F54pCTI+95bwZ0B5MoYaUdA2cOuT3ksR5tZrtlgR6oL4rEJWRbYAAMxj2I4dE
r0JEbgxbnjkvdJFkgzu6uvdek7+xu5jahbN9FKtnn5cYeWQgilLD9/WWcU0mOzMh
PK/EhJ3mhSuaTZQ+pkML9oKVVcb9RUkgGZ2UDcIzWo71+WaLA3xmhFcRdz5XMGRb
3jyR2lsXgsQEf9FNpbpMPK1pFK6AoYwkea+veJQOU3dbwaJnmAlBRJAmD323NFIT
IOAj8ZPJD13hNwH2fjO3swk3b+MopqeHt+7KbiliNJ3or9WmUxGKiZ0UiUe1Owkr
MUYNw4CE3+vNt3JKxFsVw+cqn5aZCYUudgNLXszPLVfkgQKDCQ11kfJdPGyG6EjO
14C9sWRzoYcKFZ3Z5dtyPCcFxLCTj4n+UMiUmOrfXZ6hD0myido5/atCsvr9wwWY
nNaWP4+XqUfcGDHgKum1azt8fmPATcBoDbwjqNNZuD2WVWXCrEHF6fSO+Lr6QAw5
MmH9Fvs2jZcMM67OkRV2JRt6RxN3GOwpSJ7BdvGNrdrpcQKct5pyXZpRw2YNJrCw
fz+rK7njU0Oh+ewjBZU4pG3+rvO13Rg/kdlUbx9KM/Mu4Nao4uYD1Y/17rb9tlFr
boWG5KupHcoGGT5NhHDYqIbY9D7x7i7IlGfF765I+crNFNnOHQRwzhQEgu57sXj7
U2Ugnj7pr9RhapDh2RIA6pehFZuheL/RmFGMGzHqsuhPh1JQCiycnnXeXWipbRSi
5vrxGvqHwrBj0haKDlA1M7Nmmuj+9buuBlfF6tc2C7fADQxl8QI510HDcsaMNVPx
qkq5VMqnV2S9gsSSq3DEc64Z0odMS8CHrI4PP0zSVGXpV71wz9fL4dkejXA6yW0H
DoydwnPwc7XJ/ypnvgfoeIaKUDqIo14Y/XjEfK6fWSNBMUzqVt7qspk/OHc+fKg+
rcMvKmRpBIgGmTUvSu4dLB+Ex9ZFelFQ64I67RRXrGZWEhaK0pOTER3Hwd6mDQXt
MrrQ7621Nvcc4PMaVJNZfRiQEHm1FSYt0bIhyytCQzAqagDSi11IUW666uFkSPHY
6YaIQN4f/qyiCkv9ZLOGnSgZKKCqN52AkAP3nLLYIjSfB2NGf+w87CI2l0/23al6
992X29DAs1SDtU/98iSz0X3xLOPTre3mqRLmUwL1Eue1Hm5oh8YprUsRFnR/RXs+
Is5706dRQHVKhQN6ES2QsAhqAqua2ZsqRmHd0A9JD5GlZUSd1ffU0gJ1LJrlwXW7
XQ4RmjOj/iY+7nOQgdFnaqV1IivT3J59s0mFnInXDT9AreuQbAnuUXFCSbCBPt0t
cCJVBXEaw63qUiSGukhAJBWJqj4e0sEhOME/e6itgPXf+jNY1ja7gYbs/JjnL9a9
evbgRUwmBqGW3X0NAKJH9CbB9Qtsauz3s4HZhff+TnMSVl2aMSAZavVHbHrA0CYm
3hspvJ0u3ah+jk75+iC79flwMqwg8JBPxkOTZPnfYeJg6Lh94cM07LRgGKv2CXys
DyetsPOb8DFoEeeLJL1fuRdiTe5oXlRijl7VrUDpaDo76C3D6/Kf2DCN9vA6krS5
BsGwLkXRADPrfHINoBKCEkaRWNbhrSmE+01qHDs5klCAOo9PENP0DHLuo4a92WJg
ts0fNz1cV/vGmvbAaQ4AHdo1pcDUGus7FKXty/0VCaFkN43RERCfrd60Bwm9Mzg4
IZ5AuUqqBnRwS8U1Pqq3LsQkxKGgmSke3bvUttT4ljv5nVO0sIMBSOzj8+fcyOTU
+5GclrkblNc61RaExYVfb3Nqyk5K7gkm35RqQyQdzuyCyGqHDr/truVS1HxbxjWY
/ZRjwJW1uJPPacRpMEk3eLZuKF+I3HC2Bz1DbE6L1jGfx/jASZb8e1vwRc9JOcyK
yLLbvavTHiZzhx2X0x40nPv+vTvUmIrtDvwWc/pQdNEZIQVbYpM0BP2E7zW12mwq
0AnJkWhzFITPiUTBt3qso8/AVoPeJjA+THBJ6CnQc2KMKhATUXTBAE2Orr818HNJ
roSF8jo0Sg1rdpAWBym1S8kP7umQPs+FAhCJrsvudyEMyTipmkuCk6T2z7PrRBG4
OnzcNQBQ0huYJNBPWvpGOySpCWLstMm054fQpJdT+f1JnwySq9HBTegGfyOYdQd6
jz1BJ2W6nvlg6Sy0XtCoroVBveRfo4GmMbeP9ehxaHT059rZ7oo8/Gm4zLCcaJMa
F4hiHatzdDiRIjbeLrbYy22Tu8uaCZ2rYdxLQnnnGn2FzmfO8AR7pPSq7Ah+AwkU
yXdnjc3P/azxTab2OdvhlxU3UB+aXH53klLLxK0oVBsQyiszud8AEC8MUCeGGjjI
wxm7szo38pHAePqJ7H5rGd0LuxMHsqhJ5RtLrT2pA7HtEE/CwWFdHr0ZToO2deGW
sNXLEmUwY/3czLkiEBspR8NeZxQBt3P1n5I8CgTQ39gJdDwW15vzbE45ygZQNND8
ddUOFGS7kjbaDVEZeNWp4rtc2CwhucnxniT80CgQ4osvrcjkdEZXwZxDheGNv+Ny
74gjv9hnu6GRFrfpN1hpyV2ZaC8TksAogNNUbQp6TnJBLSMH07WWxqNx26jb3TGR
JAoLRaxghzRWETLfaqXXHS8KBFiIQCjmkg2KDcWOKYAy7M2SBELq2bJWfdkvKYtq
LXibJz4oBLfx2Ppk99QzebUpzVZWrMXabPTU1cAkGBluhuS0A6tLFaN6QPwWqSwX
JkYTPNkYYhSgyGr0CVa/xNbalQMLypGwg3A8xY+tjutZZLivVQoUAj/fQU0PsK8g
u/Xy8hp8BzOt88jiTOvBDx7Zk591mziYFkIM1GWiNSmv8qbTiX1aEnJ3YY9xWFhE
sBI4CWQLk20pRfugBLPDWHYfAad/R37rMALeuypcl9uNBwzCKVoOOET+Skx3QFfg
T6ds/wvm14LhzwbiA9LYzYkPYgnxCN6pzdy/mapirL6adXsgTfGF+1JUtIuPD6qF
uDtmpwdxU8yin9VMKiLWLV4PvrRoV7EylO3pWKKCgM2usMYKAhLUBHlO9tWnyKWg
sJt2NpHRIrJXalUg4b26a2DMmj9ft6v2KboFtwv6CeXt1qLsMzSp4S+SUaHP2nxZ
nGLrH3JuNxmipB/xJIWT6G/xgJaaSUezcAUyqqD7tsyDISSaWUNsVcsOLKsyKE8h
G0PHgSvvc804o6J9lv6kY+TeY+JTWdCUDX87Jj2yJTQYOgLKAW2J85Mlsym44ivn
/LHxkZkQt/Wc3N32+ZufXNMVVSlZFvw8+Xo1ayDR0RxjXneWjYhm/0QzchL2DC7m
oPDdEJ78BenDgB6/mmZRPIaiL6+Lrc4XUuaCbPRGktlYAGn43YVA1Pu0wAufBuFp
xDX99GVaarMTntNBnyw5mgYtnExixxGy9m8Pcuxxo0fBzaGMnJ2YQdkaHdoYL1Vz
lIYfAn13tWijSMLcy7heEYW0bfVftEvp47oCQ35Mkpmap7uEPkRDuFqsvF2vrU52
NUsJVr/8MoQcsa5Tw+aWU2+a6iicQgOl0ZBrAarMmNM9rJdJjHyugARWkv2pZTkQ
gt4/Q/Hc1C3RpFtzyCZcnuRDkqJ+A2PpgQG/TcZmPq9jTfBdq34NReeXNGT8GKHG
QCdEgxac8Xyj45ioaYzthY0IE9nOWufOBe23PPMWBKr3po1lcmoEgaANNl/CgBeg
PXL/mUzd9Lg1BHHy4xezBZMB/b+3/KD1VVQGgDOWyFRLeYrKGd/nkVTuoeSXmNbx
AU0Z6nE+5pjmNNeJdIMAqWTLhPTbGD0ooWfYSAiSuGeFvHuhi9ElrtoNp+PzgZrr
AXSMErLawXpLVPrs2mReCoEcKMGk2OoYVZTQUSrH5l1IPpT0FX5+mv6erMKbpu1k
HKV2NWz61wGdmBEzO9IQrLhoHy3nTc6Fv0URRFGrJ7oEHAAtkOJQl4Tc8n21sB7J
oeh5Wr2wsvro7FHmpgmVKF0Li8avhWpWj1cp/rFuE0YPULkcrAhIUW1yDIKjMCnv
qHOF29otnDahzsI2pJ6QbBZ3m0j+mv/EA3nd/BRrHu8b6D76rngYX9vZaV3COj8S
MKltwNGzrsHbBzsdjojdkKTuNnxt6rQARpmWt/9EWTi5gFNOFUkQWYnjNdNrdtEO
UqJ+Grvh/86mwiJV/3bdcEyDx4hE2APVnaj/E/3neiidY99rLBjjc/4V3FSp+/8Q
W0S2OKCxKL7GFy44GznL5/spnV0auhAERy2jQSMz8fEudZuMfe9iXujIYXHpzlHG
BXz7z9nKzGq02ZBQMHYna8ge4rbIj3dNW5OdICH/+vwF4m6ZesMqhSIdQ8D8VmVE
vJvBFrLfdxQ5AOh5qXc4OupRjiwrurazsVZsU7d7Nrnyno/puNnO4hy+zz4h1tKN
B7ajTsyiE0WEQrgBACg7bQ641LKOI3LI4xYwAN+nmSwddUbBUINNoNj42t4UdaSq
JjUVBdK3eLHuRST6BEgfXPBwZz3aEysLLbupq1AZaPM3VWB8uY6X/L2xsX4/27n3
90G4G5WZBgib4tQW1453afFsUE/Akv1XRXR8ZEQ0J8DWwLA/1jcC01qsz3RhP0Wc
qMme/H9fBu6zuAXe2VZKZTLUzboyIoFi01OPAEYo2Gr7ewcPFEsovhS0wQ60yDQs
oIVdzrtRfmpuQEUsDM4JjWJrD3ekjnBBB7fHBZ/2xk/U5LKviTukxXEC7jp2BVmJ
u5aeHsJ+mu5fy7AQqtxkrPcLCQY8bXqRi+fjBmvaZvsJPKRo8FdBw4O3MdOcx44a
/us1bnJM75haXWckjWWdTleYuERkGY+1a09mrRjOVlq+pdF867SEqfLqMy/oAYHu
Z60ai4BLoOyDYw4z1sBX4oRjJaOdWjFjqFaa2kI0lcOdQVetcRzW7ye+YbXNtnS0
EURDxAmttnyvM96AjAKvwZCF6Mi6tRi3H/GkblEUDpzNewQ3iFrTjuhfo6burWEb
iTW83t9Ef8f72Di4fRhjJQ8jbvdvTwRG7QR0xno8A1HMKR2PjgskPWpxF/SZQBHR
xpgJsT/cprMbHRfjIlCHiba/86XP9KUlUs7XJUvrNcz9V7bk1aJk8wmSK6xXzaSM
LreAbkpjgE1QPYbzbkoXfzlNNRgw3tpvgOM34rTiabJPHgh5IjGlLqSSetKOeUwT
7CGi/NTZONRJBuns4xqiA4foE1HixrMjFwsQobZzAQ4VOp5xgvwMpzcCuW6/iXt+
FXTDCvIHu8x8Ib3MZjOTXIpiZAlBI4NsTDTc8cA0t/7e5XuSayn9GQsP1CUARdTL
7KvsYC5PBSDLPoSBlgrJfk0oWg6ETWmfYNjtTSzev42MP4hSMn0NMCsinfKSKDLe
a933fCcTKbti6n4U1htHuM9qc8LKiUMWg2LVL/53QRruuaqgSTV/QejWO0FTt/E/
tbY/oj8B1l9i3mYYXhIuoW8GTF/XMgCuX6ZtpJF5n3UZLNj/pJYTYZwu6GIIfV9m
IfFGYhYQxFPiVwDOzLkFXMTeR10+d7NjgZVocCeAk/IyWPnz6Q8fLu6OseNZLzd9
SAQEIZgCopwehOM5q+wPsOAWj4Mlo71Rab99nFJ2jqcTvObONO3XQxV3HbWAtSmo
ZnCX/IE9+Jhpu/AuAGQXYveWiFCxhmzunHpljHM+E+/qZiCQTRTujnPSjpHwutTi
gwodxNJgGbrw3LPWMkZDHHsPexrUKqHat/Jplr9wEfNZEIu5/AO3AvMpIjYdNL9W
bb3YJ7+EDYW/gXaMxWYTduPdteq3n0otfZy7kpbAd1qsGAySv1+L4aYs+mcXVqfl
NSEYZiHh947guJOvytwsftZvJ4Q0vMi5MvrrM36qf8M+k3PDjMctmT40tzrxr/D9
A9fidcX3eH00dv3IwVi49y8daH/OCwHfdpySXy91SxhoS8zkjIPaaoGarLs/U5sD
iGnDIs1+JN4StoxgzrhbAy4/QMDEFngXkQPuv7UPKoZTFqsdzxN0lQkFRjCPyG2B
AaSEbhwemLjCa7DiKCChG72MMgSh3sCV4ccJJgsXtkwCFe0wUcAhV3ZXEiRkexuX
t8IhOE4YzZUdGSCdvcprcgmD9I48rLR/CqKROGJ9XGHNfDS7UvdGnFtQ5fClJPT3
ggBel9F1isT5KvUK7mNouq7CV70zy27BlFcnIxdAjDyVl2A/xqiDwEon5oU00ugO
5hzU7uTgtRwYuMYOz1n2Xi1J3koKqw5O9b8PZJhP8MrDi0eqtjkagR9aTGMJUaAi
zyvEKrI7QGV/l8HtccSJsDWyzFkfovB0Fl8oOqMeHNSvSQwts3dTceBszW3bOVoR
eXV9opWXn/enoF68nycrqcJBV8VOEjC/D/7idJA2oxasv4xP3eMoBmVbB7Rw4xT7
a4fjpZ1nKPiC2mAQG66a85o+2kVwOZR34lmvInN4QMwZqi8vaZ3VMSniEmn89ppN
bbKzCYtdAB7j1aV2DdkdI+zY/jvXq2KET4hBKh/9DI3/3+fGyk7WhdEwF46KLeio
5Uu8ueGm4TBDbD9r5JOS2gnfBOIy6QtF1d3n0inU4K4+BjB5gFBUY42FmXvpakIk
Zqkx1VYnu0/Y1D/T22fg6tsc0aQs3f/x5NV9aZnYlcavTNBWOG7wjJj3MYNJC/N5
0QZW319RiArQqfYYuZxqW7OMRas+bEfPUActsrH5wIl0A450I6PZ8fjpLIjniniE
2noI2QWQGSifO9HA7rgE2IlcYhkspTyTuMqeusLbikejWKvct0u9kEv5pDvsiNGI
EdACo3b/AtBLzyMxXfHjNvzROw3i6NBg7cnxwi/FCFi6+H9v91Ft1SSBy6JN2mPM
Uet/AaUo5+ZGx8I6DkdLgiI7USonnuzcHtXEj+iQCSXhxcPSQeXSq4KyupR9CGi6
RJxlcH7/rVm0PyOFDcVaxjvP4moXp7A1X8KXS3MUQ0D/7iYl5/hjLP4NfMYOz2WA
/BmFPExq3IbfR1v4Q4XgXDfYy+1C54AWFpqxalmZ2yuMebFU/SOY7oJZLQlYe7YL
blXg/r/KP0IjtzD3IKJiL5tj5GKWx1xRNeLKspfI+qHprSFNKBXlzyeFQJWD74Z2
HBdwoivhpdImw8SSer549ZEqWd33RMLZJVoexi97iglMmcD5UdiI/HN/4f5LBtRf
Z5Zce/WHKevp8j/8q/7uPwfOsrmTxuhQLGnfp37xdcOY9zSJopQAZlJ8bfv+rD82
qtLxFsjz+qmezxRY61BQRTZQc0tYAY3ZicTEYwTm80RSr/3cB6ZZpk37curNT+tR
srRJKyiPwQZUXgYGK3HzYMpcpO656oytCVGSUkvWd+2Cu9ZManVTIVvuxpdPUQ5Y
cuaosXgq5nghWg8iNF3jpEzBizNY+SoeqEEJCMSPwvRqTRGf6CEif0UxadE3UEck
0FaWTk/FnCTUonxE4BAflIrGSf/vWwlCPkOng4k1c08P5rEp1XG6A5DCqI9/V7M2
8e5oNGQNgyDHT4Zb88AGSdNXHJkkxQ1jDUBtDMU6AZBM0+4WAeoAf5aM+xfhswOh
YLnqKKK9Ij8/VoAXyoKqyynmoUwaq8tOx7I9QznvMy+fTtluho0CyfO439esq1Rj
`protect end_protected