`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1456 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
2mA4eiZXfChkavClTs5gUZQWlsEFY+L0D7i6MzWpMqp17cfA+D9l2u5t6PjAJpMb
K7zVQCsTNl3uFXmFWoO6yGCZphM3stdYPTcNDxyVSlwQvqqIo9g3w0Rx0VyJVFzd
4a6Wh4CReOjdnHk1pOkfYWxq+laG3q4/XhWFiSkfYnEPXYqsBElUUycWRsm4H1zO
jzAptS4LN4PhznBoQM4y9/sFszncZhNmU/CZY2TvtW85ulZumuPCMWzHFa1Tcdns
l1/LqmVWCxb6tvuIwz69oc7TT415A3cmInB4lkUdaP+wjbVG7LJ6RX3p759zTBen
Ah4+1ikSiLVWPWykUJDB0b1rPbCAm9QzTojnoFGFNG8M4NccyeuSQ5vlHuQScDKV
5Hipgo2OaA8ald0wG3Ue6C4pdCdcJ+kA4SgV8qgTaSpBa2NTkNjDdfklpLG9Tz8/
7EHJQiCZ4h1N3nHhtsbNvHIdfVh/x1mFZEdVkwyukzusm48P6mE7a/zES5ns1q/h
MfmzrgzfnTP341YRuA0QuAxL+0CEe+9Vvkne5UAq+qehfkl01E18Xpylu5SEMXfd
BceNTl3jzY47IRwFjkEqX1zD6+Rrjm0HBgcRKysFQUd009+K6dbKJy5wycLp/3cQ
1JHojGK1/xd/F6GpVsAvg6Gh7DqdX1CcBm7aJml7KSSmvESMsXe7uS4OqPzOCGBw
cTGCWdFa9Ia5vhs2zle7WTvtTHMUkFkvQ8iGQFVYXea6V+SR6GpIGAEgLTquyXgF
w17K3OTRggEQQu4fzIEMmASE9p/vlUz+TDEI0+WkLJR7OOYp4cwIcUHCOo8yD2a7
z7PDac3HO1jhlha5eXbNxIOdOuNm6f1Eo+vj3ievkhdWiTilDkS2yW967bVEJLjq
fiCACuphFXYrCn8EvyS+0CQij3YF2d78qT6V1fdJ+z8ZaQzMda//86/dIFcp5cML
k8NvCJ+lIF59Ez5fMQn/5Mb04gW/MQuHjHJd3dQPeLz45YmQ0Ey815AjAqQQRRTY
aTWhs2Bdly7O6lotjyBk+MYVq4xwT9UbTLylSWxQ9MlGO1Q3SnvV92DhhYZ9buZ6
qAKhBMhSkwLd5xJLB5H0neKFB/shScqAxfjWfAjlK3ByzVmQZIYjitLfh2CzpgOJ
R0n8olGk78YMRFHgi7gyjY4gFPFVBFLQeIODU7Oer0oHZVTcxONGqaf7/DZg3YOl
QEcTe/43oZ0sFHtgsTCsNtgCR1ozk3ae5BHVAS9aaTDpAPqcwBF6VZbH/srOVlno
DoZe3+DwA21vhZGiNZK6ijgKdpZ9Vqss+LID96dh2pKeLGbNSSn5jXEJxJqj9nsf
qzc2z/v3owaDqvwa9rtHBLvqlQkuZZGmeudxDclxP6axIhY2+NO3uaY4H3h5UseZ
ZMKLoeqR+h6+9DTYpwzezEYonW6gIzQrPBJFNqL9WbDKzDBljX9U2jDEELmbTdjW
5Q8hoHoHHuHbEha88CFcURxe1GjL3asH9JU5avYLCfgcGsf6XUM4tbl6p8LZ7Y2E
MgM8fGvazf5uO1xeH6CDVIXCVNOFgXVJ5bLbF0+oKxNGlZcg6SScQOSpitM0CiUR
CVYlQI+MzEzoMODTqr6UbvLi0vAA0G18Sc/SHfRbvpWsUoJRMzosrRncB0Y68tsO
jJ3ECquZ4EeXvUuek178cI/VHvQpctmWGAkWlPiybGukNqXBwDOGgAN3fz/CiMcQ
2O7E6vhkTT709ffav11TJLWjorbG57pybK2FaORRS+aYmpcbV5ZxSAPRbvkDzReB
JSHpF3z6m++tzJxMXET9cA==
`protect end_protected