`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4752 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eislOGByxcl/gRn8UziAa+H
mjgbsd36EQO5Ail/O6Xu+Xx/ROMSlvuBazdeHDaf8f7V3IZqPZclnVuOx7MJH9IN
owXBqHkZpMhuah7CAFoFGbWW3+Gg7vcv07JISBBuzCW+CMjMTkc+XIdi9x9OFHj2
BAaHWDNqBBgVi/cppGWqxD5QO/rvwY1v3M6xSQ2DmvADJgCFsQT1ErsVnKjLul0A
CIUyQft1B1ypi9jMkMVVjVrgGgUJxAtxFWseI3asq/0UN6Vbrtx97TXNUXRYn6Z3
kv2vWvSMdJQE/M67oTsbcSP21QHaoP1MW+fWeK4S/18XlOyjuJf2z8CLG8A1aZhe
SxgQjdXMXZ9/T2Chy3rq9ZLMpsaQA2kVXoQIqLwRiyVDkTxjDjOpmcvQwEFaKu60
KObtdmmpIzuqKmmUrLgO/LtZomQkkLMWGbxpWnkE6dYzwTMiFDSF+7ms7iFFAA/w
h8xO9BaQjksghRIxkmjF8xwvnW4LbYjNGLK1E8avFStBrnAWgH1QtJcG2wAKlp0F
jEbGw3w1cqBuvQVsyfF+HvAYNbOT444wTTc9n/1q4Tf25bWe3qGbFZLLeheq7ID0
z0hE7iKjj+H46im1EEuXDRtmNFTNEFDc/SVRZ0ZO1kpDeah/hfc8fcqPlH3Xgjxv
QNJKU1/GlAYlFcpdTrQShNKvdtlSJ4otn6q+AVMOIKBMxrFPvnt8trXAcnXPwyZW
PuFHgu86vC2kWUnFTQ0LB9le9JYPKqfaWV4AIc1csy1s0/9DXtG/gkxzKdKqGyTV
sXe++Ci7udR95VmXuDe9KPzN01CddlwRnGVM4lZwstjR0TxYRQ3y4ru6GVDtNiAY
3ujQsqkd74uldoPCDYf64RZ7NJWDxgFtjA5zdwJ6so6eRE5BEGiwschO6K02T67r
wJyzTB9Cak/gCv9tvcLi1UiHJkaVIF4YFyDdYzsYwW1pkgc4pfViXxPsJa0s2ZFQ
9SPTePNoJNgSoWBl6kZEZF1nnKWGHWT0YlLx+nxvAaGtjS3p1Sdts50kel42VeGP
FnkqZFo8Ue/PzUTAPwGhlElfAr53bN+s3OYZtx71KxQKNZyZVpB4n9U2ADmtyjOi
F9Jo4eU9a0vmg9XHM5x3EShBNhIv57ClcZPA9bjVGtq/nKfD6ppccHpwiA9TZg6U
c/xGoBCH1JPWpqn/dM+7vJfI1vmS8RmoZb0RQjtFszb2Alr82ymWAV2r09NxbHga
L/ka28hEH0iSWtePUVz28NM8lCBH8MTMYTOjCTz6C9hBrTaRHGxTe9LTRUkkRFdR
M1zT1w9tXGgCMIaa27rfHt9o5mORAqIGqF1W9QcdCxcPQTmf2Q96SWvsO2ybYr7Q
YDJhX4IP9qNH2tOX2FJlmjJciLKrxYJK6wAJlP/3I7VtPythp3IPdstdwLdOn6bz
Yk9J4NejmzfacrXhOsEbJ6K8JF99094btQvcFCxxrxkTwjHqe2QsFERjjnvivyIU
pkVfDRO0twh2zNRZ/DKrL0MCvejiz9nsIE4cuynjQbE/Y6D1PeQ1h7Wvt7pT8BHJ
DBVsZJDzMqusSDN23As0iqxe2j+dXkGciMYp/JtlCc1nhICdE17sRG4VLdFnF+aq
5/mP6pU3HUEzas0luZegjaCUJ6oyzs9+G+KoirU4EfBidmV12fFYJN2xPztOcU5J
BRqEEH4h2uozQh8a4BXDgr0IW63Ps3GKu7PSwFTprtmGC+27UE0bi7oUF2nAobnB
yMia8K6jfmAGRdRhi1c517mQQHmfpIDzswWR5sNA+rPlpms7Wk1nYHeMtIjRFE1h
7aWWA3B/eooXFoDpd4TE/AQpLwfIe2KAiTkautQpSj9nW8YxRSAy3ysnKV2rK0FG
hWdBK7QHzUNWOIpSO2kXZUfHr55sK8WbZVD1BbKw3zI5iTUyKGXnQyCI28537tAp
DGZNWxuZxGsIzdE4bLScW09te6Rqigh8DdcXe2WNWbhHFx9EKkfdI9JGBRKFgPd3
IM85rieCx5jMCj0vi6jRQ9Q4Ci+g1O6G4HV09tL6nimulBlYoM0jGxLimM513CPn
p/9R5znsmYPONLErzE2R6hQThfE1L8hgWy7hJEQFzTjuP1T+Q74MWLLNzQvyY61V
xcojmjCtyxIgxruBv/7jRQKZlIpMZKyZT5mmy18K36SIFaGzF07l9B5ZgqdPjVF/
KpGBh463pPvie8VoVtBSGn7y042bVu+cHFdGe2pWGheoO3n21KzysIsami/+quxj
MeIHIUUhjJ/GD3//Yh2NwoGYjWp56r1NiQSdT8MJmSMXdLIFl/mpC2Z3ZAWISHTa
vG95eW6uJ1Vx6K6z8EKKnoiUQeJ6+ah3RStFq0+4awzKvLqIYX0NxGCbdEJ8uHF5
SyTHnQGyWmfgZLCa9vHlQYbjDOYtmr7gPJ7376A7uhL/y8L/womhFpSu5xNJNyes
sWIWMw1HgBa+7x1syjstD2VQ9OB9/u+tZBqxkqMH/kq8158ZWJWi5Ur7HcBzAhUo
KrURlN9aHjnt8yrJL2BXV1ZT4boWdCX8TnMKDp6lM0eMsrmvi1eTkJK8H+yFO/Uc
Ag7msPGx7/LDn+CRiNRt59ekw0n+Pku+uJBLz4mYPH0Xb8YrY5iuIqzqFNPalxYr
2+wcC3mCJxd13F2GENNILhoyFWMeWuzwuq2OvRtztMtochdkNTua5gDqtU/US9kv
iXSnVwdqOpUuOChlJEQVaTnQ0X76xyIyxVIlI3HtOrUIi5Lzn/hNn1qT5HFjgaq+
EF5g6boKnP1nttWwd0cRwnlodDcPzJM4RTkyrzSPh+o0gq9h9EoRE70N8YnMOveF
AMOYJFv0Zcxx/Wkt3Si0U53DzvF8DsEbwksaG3a9YGVmdoYQW7Nf0EkJHCAu9WMV
G1ev7dazMfbJE0ugJZtTRf8FWZkuNIT4Nwc2QKOQ6tQxnxHbhtkkP1n0lNG2zTh3
Er4GZjX66NCyxUZTcYfM/gDrJd8BcT8sa7SX9hr6o3ydDjJoSyf9K836suigNqJP
1VUOSapB4vSL1qP+4tmeaCaYlsZwKfLvnW7DG5K1fX1F80jeHlU03X1x8js3r5kI
kqhRVeqDMOCU4Px3VWjCZCXmWV7cpvmvpBcfXSgAMWSi5Zp2+GsTR/W+KoZyxa5J
d9OYn4nIFwOrlZJ1/dQ0oSIgS3u+wyb449LX3mAaeG0aBcLKL1MNnr3L0n6bT8in
Yy/5wRklbsHxL0j+65MhZ6yX2aQlU7+i42gVInw2TlA/YQtkXRAQRQ5d9tDmcRq6
qzkt4M+UmkIcDy2MIWwy7OBzLmwwny4Wvr23cdogi/7/0pasBGJDRkvgeJVhClm5
R+suDWVssAD6Ckb3L7SfSK+/NvHTQ8FKyZRndnyLq1fIedkpvNB+VuQW+obiZr7Z
PIgdBfJwUe9nbL2Y7DJ0dgM4Cuf0z5Z5xANVnzQ/DGf2ENAEsINMmhOC/Sw08wBY
1yPs53TYgM17TWER7gfO8Ec+e7arhhdZU7wsVNPR9fZaKUDRFJTIzRIM5rmW18yi
pT0J6jFXJLq2ym0ZgCz3n3H5g34k6pbZnK3C+Kaq2sI8VIqVYmxd15kCC+dhk4s0
nsU0rIEGRf4NQxw7aK9kLfCrXv2hR4R0LNAcF5kV3xfG4VrzRo+iFN/YIunI+mqT
Yz1gFsDhQsWRwrd14IX1ilSQAvYrabazEKNU+Xs5rk3AVE9ssudpUDy1loMHewwT
KnMIivn1uzgzt607g672FG3xAuosXvS7Xgl6+AQSGRafgVQWRkHmBQWoSEJjxiaL
itSVCsasLCBZznyaNdda1j+3LBTTmYf0NgtNfT9FhmJTzmdiTxnRZ2XUKavJ3X6h
8jsiRKzj0dlOqx6vBkml9lxIt1gFMvQBg4P1bPg3/hbu5nXM/5ZovUADMI1L3+TV
RXqsfFDpARS/GE0Y0+LEO4pDwIct9FzUNm54J858NvjL2oytMO7OOE5Aim3+IzWN
TpQC2idNc+ZfgvoxQfsysvKcBE0+Ere0oKxdu48PKtvn1qv3Lo0Im5fDrcjqf9b1
L6DbpjeLd+tnLoOVC5c55mutBikqHBLpRYBiDLSHGTF8LR6XFRGSffQ1Lyd+vWYt
N+b5C0Ye3bARge7KdfO1SjKaZwlUirjfH47cGJz5kmmslJD3Za+h8wJUYq2m1w+C
BYGJk8GRa98IVTkMRK7KuXedsG6npVo8rYOvgnzc+jfRtqjj2HQGrVSiOCyy70G1
nfNFKh2aCE+mHU2R62UgbTseUY/sPttqLkSuAV//GRfnWkYlSWOakgXvxb/4eQzh
nWGaCYeI1cvAwQfbLkAlJnhssb97Vg4HerigUiJvNjCSQu3kke3zBt+OGtiUlnr6
0EBI8/dEAQofvpU68amBx9bof332Ep5k+wgIn3esTEuOhMQVm9MHUbKt0h4ZVMA5
mciWGFFoJ4U3JPZFb8yR0jhXBbJSsTSpUUj2oiGqt/6OuZRlrbsLL2G89M98HMrb
TTby0vnyA4SJOiJZElXNwjKi6daUdmtvrLAKz2Il9MCkxdf2HXC2kcn8d4H1ea5Z
riIA8VK71oArt57xdYlWiBZ+ktw8D+9B4E7XhmBznOpNVHyumVeWuGWLkyEbKqFx
PJ0/rHjM1oWoDQ/yAvvl45mf5qUKKMH+jBr4ML8T8oGtxG1ZWEZuvfbC2pdY6oOp
ss81BnGxdqXp/c+2H3v8SEsslQnP/cZhb0L3NOKE6X3fPEAAzBlr60q5sAp6Xqx3
16/B3bll/MeErnlJrAZlAVzf/B3b3/pJ9WNFW+QImYI9DOlGR0+jjtY324De97dB
p7i/yf1x6sLWaSKEake3GP+nn11GXs8CEjEgy8Bp6lEOqVAkIIIcnFu1ImXa91nS
9ANZe55C4TIW7upUFdj7fvs+taAPKRSmh9sqVTosPaxOdu0b6gTM/8ILKsgo57G9
/ZWzK55QY81Xvt1q2LvW80yNP+0icvVVjq+fQoyE3eoXdIr5ZQ414pxpu1ETHqlU
F9G10M6cZpE2IQ9SiyNHPBe5ovqi6C4GByvQ6An/KHk69Khj6FM0DtMxv8Ro914D
PAoE/BoEPd3b0GP0mQLnni3VaQ0GfTIKBWcjLbu0buD0UWCmiTjOaRYGknYTAv0o
nFlOCF4eZsTjhuFryt/SNVMO6AG8ns6ld085muwOP4mPgYLOlBC6p5Pj3zt7yWwy
M3uVcD5nqlbRmGLtOmxbG49G+wcw0hveyWWjgWStjCoRafoUewm417xHNCRsI54u
wA7tKtPOmEH08UmozmC14x6O91zRn14XI1n+uUtKv5uaQ6/NgTEG7NYvzeBB2cLQ
PZP2pLbB92jrLQoXUqnKdNcsYXDSXyzcSDavr0FJ4b9n6lIc6fcWt0ihj19xqIeI
2huU/iPU3GUYlmo4Gwo3uyW1j2imAwHwRBLJuLO8Bjv5F7CZEQQKZXy58FUAVfDI
7lCAk4nD6y6cTyap5WRhY7DvoVYIhSZeTw6SXWJBc+pb8xJGCT7LWHYU2Iaj5slm
z9g4Fgsk2BTz92p/0qMpdxZhNQY68z8h3JmAIuWjWkZnYqtups5DlT5gkEhCHDAl
8Hb6sVqSlSn/QwYWZ4RUrlypV8DEov1/1QjBmmXyNk2Re2RINK78SIowXhJuISie
n93+GPLZ0yKieB2hOdD9rjI8pwXW5aB5QHBtdWSuf23OMDVdMMR8efsgJibIbjvI
VJ8vQeecPRKGnYkpMnNHzmohuYCiwoIBA3lCJXyUKiivGUEfTZptN/+eYd5XhBOs
l2UeCsAIPYv0Oe4IE90AD4TcoO5/EGxMLymtGWcvmpV9yeEO0m5ti1OmVWhYfkD/
ts4VLvNYYI1qjSSIMeKWFpRlOzvRszhCMf5WkOH0KLlUQi37j3PbyG7LQ97iFxOA
5gdkIc+x67aUUDV3SjiIcG/ve6RvZvX0Ib1LUrUyoq0CUtFQZXMOg1WnLzVd1yDj
QwI41A5S0iBGyXxtEXKIRtQywd5HHA4y0+Qa52h9Gvv7fZKMNLyEUdQkXnZH26TS
N3x4N7EDy9VfPkunD+yyMFFOFE3VMaHg2ugwosZXgOAI5YHbAUbo3XG3JklkNYTd
gQL8RAhXHED0IfaSsMkXYtLp06BpFt+4yKqCogbtpbMRDgtoD3rO11HclupfgbjC
bvHDNsrtUX4/2LiPv7lxBxh/GfT+V9KoJm42IZh2woIlnFj8MXR0WsvOJI/Y1IfA
`protect end_protected