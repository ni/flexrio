`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 10128 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
S993bpJjwxtMDn0RNN54XzRqn8HeK8t/Cy1jDqZNdl0d2Cg9JE9dxx4gcxgrs1bH
u9okuHrVAW9bwwe+KNbXSScRMf4Qm9xESduV6RVTlidG1IdSSZEFJfD7IZqURrmO
SstAkqNE0j0UoKihnCuMNItjFDj+lzBOc1Sy0D4BUOiJIo4SbPUnU0V9E2+nFsSr
4ZuxljlORVh9eluy6Ut651QHxw/Z+9f5NTYo3tjyHd/EVlALriRF4yRO/WVKkzzQ
4h5iQolPz4DvWVgLYE6w9vYP7U7dBaopBh9YRQ4/O9xzupGqZRkVKSe5S24Yo+OY
RRn5F9tO45m8DPI7Fp+9oh5DSqcABk381stG42orv3BOe/hMqT1GRDOnDhXzcMyu
8Zeind85QfNvNbsxBMRmrapHnSwj12G5fFsIn2MBi2lpVg5QvL2OWMOTInmUKJtp
m526+N3pNI1DF6k2li4eEBf9mqrjl6lSUoyPU7WrqCzPU+uOz7TvmcyARTUegGK2
q/U7L1kd5kKMdFEsBC0l+TEQ5d167rQ3F5cLR3DOpQoAXfF1x9Zn1UGAB63BiYDA
qJuVN+WrwGlKrpNyFVX5+/JxuFZRgGlgKGKIIOM1FzuGi/o/W8EOpFN6/B6piVcg
fHLNIeCoSd5POYtw0jNskkETqOgPhzhGxeikw9S1CgABwS64owYwLqe67PYZPU4V
/nzskjTh3PiJ9gbPUYE7Cqk3vtUtQ4mKJInn7xTL8bM1zeSCdUz+QmKGhvIWrPM4
HkKxAH4RoLCkYiVCYBVm+WuNrKA4xPNQo3IpNsnpoVj7KxWo2wfMEsSYUGrgSvcz
64tADlDdYaqbbTQaD6IzWxKPaFhugoz5pDoHqiKRg+8jdXvebaKmQ8vnGkN12yzS
kILpHd1dorlKHfuuBDVP4IxosuJs08dJOYPoUH2pHP3l+LwToPKP9Rl2ASLsqbvR
HfOL6WEKMFQt0i+F65vX+MSZL4ByYS3Oy0+MdoOmfHL81OMcmcINGHuitDtigPRH
o+vE6rbvUzyYrZu7M/AC7Nz+WAN4F2TNXWRozz7MQcmTGIvSUXfeCbBsQ8OPjdI9
wpLDJiWiBDpVkJk2PYBpm9AuQ8KnNcTouqmf4skA31B1Ak4IE7x0vHmpvEke6AyB
ftyTBsOOTwbepWYBKJkBViv3XQ5xiDNpjwcV3vSwSMhWUbuC65I5MVMIMnTnFvds
f8RLbd1XyRn7xTjl5BFDIrt6C7OPUvOU2kPvG3up9iPyKXk4DG/rCF7m98Sq8e8o
AW0H63pDV7t/SuEwOXn28pInNOH+dVHANyW2NspOaum2UskoKsw8eGpeCAll6HWY
Rmp9z+8pHmouvePalIwDjB80Ki6EAKf/+U/jnS97zmn99TwI684xfauDIL2hqwA8
Z/AnOzxuFZlmdpew0Rqv7mpnY34TbCRoFSAguWEs812oUabJSleipPb8CAtnKzne
wq0gf5j8xgsUiDe+srBIZeciHpkro+MNKv5gFjEnR5YneX/srtFpjWRx6JTPnwWZ
Tm4WKTGmQh/pglR4kuoJJxSp4R8zwVpOYY/NjwrZ7EYloRfmEhXTRVmoW5suNnuO
Y/qO9h5cSGX6osAuyFmOYD51kfxbz7F3zXGKQFQlMCTZ8xR/awca0UTCrYZELWcj
3bdPq0QggP20GqQRpKXr17J51o3+iFDdA0w6GYhVAuQTf6ACv40ty2Kxartod3ca
7sWMnnHFjyPVvNZUiSNca97Gnz6jr82zTtkLdRc4yGkZXcWliGt1mYJGav+z2BiR
NbCmIypHv0OUk0tVkb8CNqwR4eAkymzGdYOOkNyv0U3k+gutf8ln2SU2qZQP0mIz
3xdNPsvE9Gan10Bwc2RbmiHgj30NxgtzqbiS9d0FMXhlNvZsvh1RJQypY93/0OlR
elevPpMjUt71zRIgHB+QaffFTsi9ES5/pw+YqI286AegvaEV2vm8/np3N1qdfAuU
yroJm4jFRD02eXogi0HnVe8IIwuq1jNqDfuNtKuNJa6pkS1Ct2bDCf4OVKLukG1w
U2pfqcnhiIxQq4q8JRXUkM+622Q9Of/FMsHFKW0xT5TwgyxCCgi3XS3l3ig/Y3X/
Tvjl/Yxb46YrSuWRX9tpD2g64PKNegKDW8VEP9TNmqZsbxDiSVaL1m3QcLRs/SPe
n3I64fMO4XWzFk9Q6kfv93b7p9TgSyLWz0MhmL44VARL+3jgS/wfO6tn3/AWkr6/
4LUYVVKB1SJKLdorV+ttkDCCTJm+gLyjBDU8sZ8phfXtOtA7LqtvfVZCSJFtU+Oe
KrBVugxDYSXIdBs/Vgf8IAjjB3yjveVYUFYNnX51GRumUcfrSPhhLIEh8f1Qe1/e
LtNx6UFrUI3gA1g61h/HmFTAudEfSMuAL+Ug/E2pKOYL36O/QzmW9XCgvYWUQhbS
WHwp4U1+nlrH906IcBWyXo9fcGw0rSzSal8LL3W8lgrlK/gOLefeVEW86R1cOfY8
sEnRFBPcF5zK3eOVQeNsIOkUcrnCwLcp9SdalEV3O4SAbcdErl4FHkfA1LugLalH
W7H4l5HUVYjUkZ/nQwOib5kx1yNW7+4iqytLvRG/halMU+/o+76OjbBrgAPOPGk2
SwqpXtzrXtlCWcby0pgVaCf0sc/nZEPsRLQOCfcKyYdBNWbJYjTDcOfogxojd2Nh
73UZPPC0ivlyb+TxwkHl92vjA6PADyfKh7/bDBt+/9EpJ6aB9yUExdsFoQJ342YP
ekWXI4ldQBb6pHY3GR/7AUuqgKof2326fCnQ7r7+l+NovxMIX3St+ss+d0XvlTA6
PWY+7VWmG81U1UpBKLQigbhvNtMXGZXyp+NNdENUWPgriux6BsVg48ZRxoIvuow5
+xT2fSYJQOYNHswG/IS0gBuVgkfVtNqVJUW3m5NNzuP+LqQDbRwrz0dDefbnlJng
TLkISzARue24NpVCSqlGHFT1G5eI6fUSzpmeEKCpjUOKIfkYygpyzaz3sXzIPQrl
BQbDa7w2D6QCw3Uy2JjPSmePpcfK9LWCnrdt5oauTHlPeiMzGCizEuHp/U7sNuHZ
sw/D8Ux8x/f6o8BgRiEyfY34qcjk0/XOaXGEZXVNeIPF/XTyDhcRY+L3lt3pp0lE
n1jYqgFujeVhYhNk02rhj6t8YVUyyZ0RZOR0kiCEbm5tQWlMVQaycmF8I77VyRbm
sHhJzkTCUfVZmVrq8Z0TXotqlvXdYAIxBN5VaEjMQDVQBZq5kMsop21Aa46hVZZ9
U/IDbVB+K/3FUQkjPzSsqWmj2SwsJ0AGmd5Db2JjSAcdUyaA4BUOrlaCbZTog0pc
4vttTB6ST8uE7Pooc38HnxivHnsAOEbh4vYFIt2IFqkxAk1wACXYgD3sbY+3Dxyg
Oa6iwlRBc3OMCNdQeBbZhMiocdD8Mg6EWyWd05Wglc8/vozHgfyaI6Md756oaq64
EXx2Aa5bwAodH7NVVG6v+0VBi8u/UerIKGSXUHA3p0H5RuYHGJR9HFr9j23KmMfA
alS3Hc4we7GU2thbKAtkzTMCbhicAV1QwyiA9rPF+h+gxCf3JtCKA4bKOgkp9/WM
as2YQ9OahXH1PoCJSSIjgdeXMbvUNSzgBuqL2zeqwFCOvLfz9pdKO0R9jItRg1xH
Gv0eeCYZLM1t2mQ0biJuS95lqWHlSIbZo/XO76QuEOrZgq/H3fTRYtKtLvCinL7i
jJ1z9SrIGbq/Y09uRjaMPCm4l52/Mmln7OAk8fm7vxJAL1c3I1O9pIyNVfEe5pbM
wcrv9UqgSjsssPYJOWzrLj2jlN4cLeFlysPb+v9BJxp4D8W2LIxqG5ZdOL9hJlUW
jX6nxC87OtHnGn6PrlEL2Up/jLL7Atv/slHriYbVDIo7eeOqvYYPjyYx4sc4B3PS
v4tAm3Ncgw8SR1+l5tre45npdNLadrBowvmea5dJVr9GtalkhxYgFZ9WkSszv9YW
tU7OyUmX1/fy8R5KC9tV0laY1g788AIqDD37vP8lBWJNVvh/tt1M1agc25xCkI2l
EAjmp+0KpZApV+KrQZUxkfpgSENTqqH0rstWa1uiNRioCX4wNB1QDIKyL+Lo/0d1
m0dtvo0IicCweh34YlT8zWHnb5bWE7lc+0/IbM9yp2bWC2JUzMEcN+/iYd+ZYUPu
SG/E5KAUQxANqd9VT/TNakt3C8Yr6wwK3ol8gPF1OiOS56fBXG8GSfU3+e9OalNE
JPZ3NAX0RCh1hL2jpcX+5OwH7tEL7vlqB9nCCWFlSoIA4jhFHnwQ3TVb3kYMWiND
h5TILMUa0DcARnLjqONWrCPrNbJvvx2lktXS7upCv42e9pVzCl8EfV+BDU+ef0il
CrMyvTZt+5fuc8ENhfv+eYynlWRsQEfU49SCw0df4RVOTEA2cy3bZN9ByB6NrDXv
kiTE2FFC2a23BQhh1a79EC7HXsodKsu6/Od588bQe3gaRnPLP3bah9HJ5iaNUGa8
MNzTdZQpbiA13jVtQ6k52F0wXvp8OW5BZV5lTGyBiyc0X/hvfh67FrjhnfHZ01mR
WIIEZZM4Q9aGKF2xY6l3q0dsjNtySbZ/El96YmwF2ywwU5NmBMUB7ZsY3GNzVrNZ
Yd/wV66LJJg0LTAOlxkk3+EWsq3ssOj/SgO96zsOXCQBzuMQxTOMpo6iGmT+sUg5
ISDS+EOKaB9m3ENQI06Jx48uUwv8BBW4kl91sCPbgsG9iwHWEWvgar61HPmfqpGZ
ryk81f7qg+WcJG3AZ14sjI3OtduZ/ckvH9ICy8FPpQOTSvAFN0inhUtQm+QzSR3I
O23E1CjeJypr0Tdgs5Di7L69K+vN38P7hOBjyg8U1WUkdIIu+BibZEkgRwbpUmcl
uop/vbz4daxcqWznBGdrUXb2G+NB92VLoW9FOQ2z21iuUHVknFahy4fgV9bRz57q
4kp26tp2ibDESrCwlekRLtctnEu7RJoWsjjhoe6CO8Lp5S3V6OJashE1IX69Brp/
9UCsZrNrjGQT1GOtygR+ijmOQM7Jh9hYU0nCa/XjeH/Lz02dhwogQA1QGpGksFUf
jtNoJUmlYv8OThloDW9PX/w/tNTaEWh4bvVxCZv1F+4dBqsDq/uTpXzQdjwCEib7
+p4I5CdOqMlyi/6GHXvXzxJMeLZTkz7nYI37klffmRfXqEa2ItyoYEaScWs4P3ay
apRJ9tu38y4nFbOxB4PrHPRDESJ3d+G3GiVbPKEyJSfW6fZy/s0otVmiWu011n86
jw90s6sNK0/jTOdtYA80O1z7zZygMfbwZaHGheTOgJe3ugi8FHHcZ2L8FoX+CzPC
DfsZQ0h40E5W04QFZt5H/wXV7h3JERHAfKfdTVdTZFnwJV8CmR1a9KBFO/TQwXKg
tPrftusd+ggmdsFyx+OklOaARI3ebLp8sCQqvmHsn7FQw8bYdDPOIwLY1mYwAvYA
0Zo64rRReQ313rZrNJGBICbrAshFTCZUmqB5lNo7je5TJz7AbOzJnIWOBgWdHpRm
17NLZGRd8IscbATFVf26sLibes8WGR00+8MGf+ai+mzYK0nFTcMBEgBu9NUtD76M
rabj5J+R5cu+EzjClEs4Yp90AsX0oBM+MSnflNjJ30AJjEwQ8mByp/STpINWms7e
6xf9pykkor6nbv3ux3xyAIF+I4MbxfWEarRzbL2Q0O3g+ztgLt1JlhO6B2SMct2h
iCQ4eSgkzqgVmscaO38N/yZK4sEXJ9MyBLKeaIGr8p0xELwT+KmArTs9Ie86IBw8
y3sFJ1h12KIGCuiV2oEwvc9dHgySL5ZDxTZv6rR68KBTDJ6cLCtxVuJ+84eAZ37x
VhkDdRpuWFkwDucNmh+KBJZDbsXVfedWjcQGLzCj7oX7cKcmlzd2pRtJPW8lPVzH
F8hWBWZHV6IxZCJBg/ai8scupmp/k0J6ZTD/O4rncVR4Sv9zuwvxPbEDlUVL/N/4
/GVMwaV1TYry4QX2X02YBxJeM09n/ajiPA7HK289tr9T+Uu+2FUjo16SmOm8pG83
nglcFw/sgwZ3yaxTe8flIZkPIwiie1X7W2Shzy9IrUQFLlfHGZBf179wkYtZIDrM
cn7WNQHbACiPYLEIxAqOZmRjpwA8NxQV7NBY1p0MGh487PmEPI4+Bvy/57Xvo/H/
1jbGmuENMLsIRxxa68m+Hi+2bKzcl3S2/CjQmEpFV256CukjhTP1oYlq1laTopj3
oZxHGlB4D+ULWvX6Bx0d58UA24aiK2l55EUNM490PKiS819BWqB+mZ8/B7UMtJYC
rl7b1vP8v1Mzt97QL7nSXSMdj3CgSZ+NDoOGrZNtKigv6TqtWZ+srhs0uWjR+xoX
gGH/LgbvDU7NMSQoi7zJvpCne93NFWoAeMhb/UEPOn5AOCWoT2iNhyZRrf+ajQma
G/0zbqc/JC/9XWUeKq84o+Gf9muH1CVFdWrVZhkiP6H3DywNa8XMn1jUGw+hoLJL
X5WVtA4+aFGFu/3kqgolok+fCFcrkBhqLlfg+Y6LutmWfFi1VFBz9ab46ce8bcNX
CGX9ZLcy2LA2oDe07oeACsjYNH2PCaA/E6Fd2Iza1193UcoENsY2b5U1bF/BuUqd
HSWD5U6Sw27/nqk2YElTAyNDCY6IsKvZL3qBptFDWK9zE0jWyrL0jcnmC1F6FmoF
12gzoDoEIDVdjVoEPTUSSAjR4A20hW2+bIwTT/5OyhSo1UtgyJx+9lWY9vYYredX
rudZC7ZaNo7u7UOkyCouvQ+VQCOpES4FQ1epSHZnRhna/ykq6H27G/TQEhU8rIod
mRdaVG2avKNnG35C3lf5RUj+6O1M1m2OD5iVUSULTKLFeEuTbuXKuE0J/jqtKN2p
lDeUeKhrLLlYF3pV2TDIuUUcwKxLk/viNzKRUhyf+CVeq7+fqC9jgsa1ljZjMon6
e9yi+UURT1K2zTUZWv1SrPa/9EFW3O7pDLxXnwOEPGmNTzw4V90xC1KcLShvLqFw
4GyouOls/gsz2umUaZLQPsOtddU5Yzd/zcgbQhUEd9bJV7NpXgQY2TNDP+xM1Vxr
wla0w8fPqlcpLHsARocw1zbciLhZRsES3sxzdz0NnDPub6VLA+7r874C0zxp1PT3
tA5u+EeprrNNTrjFifD61vHL6boGPnegDoOBuOl9ydqHWX4RnRAAGBoUWcmoxp7j
nRDVAp8ButmBQVbLnRsMr00oD6esygwcvyDb1fF8vBG067fgs8QxJBv43w6OY/O2
RUPYas0uoScqYcw9IkmvTkYgIp4yDCfOGYoR/Hdj36BNJwy3ZwI5zu1hm+2xSVvl
71S7ERh6SdPJYNj6zSTHVXcDPxWtDZHD6JEGix5ptCJ0gOhD1m3Li4IEioSx1/dv
OJIFXt+ctXzgoYrKivz7sVUXPxr1TaqbeSXn1YcaxNj6p/YUKdyrfZzWpGHu4169
PFrvlJvm0Q2LDrx1kmlQHMKp+arewJRBNKloQPsTAdMJlb/SPVk3+tdbdTJYDVLl
00mnvVGYtiRgZe/dPHc0tFDwx2gQCS21ePb+7o+YCE9QaugQ7V6HfxfA1KgUr5KN
5XmhvF2r+WYX5MnTvGARspzumC1/OZESLJgVSOvtSuKuWHkW1EE2BMohGMAHI74O
Q6WVMGEiUfdE9fOGO0tBcHbbr5/IrrAoZITzCdE+bVSId8sNxCu9gKr/rPye27Xt
T7z2GApMuWVFby7eJm2lJ+EvYBGVnEe4nVI8ykTuwlPAhApu6Z8XBW5LZWG8cPtS
3iHGYNlGKVV7lsPlG0HT5uiiMITWUn8zXmBAQmJQD1hqT7h+EOCt4IfyqQ+YSE3j
ZeL4NlZMZRhwowPXMjTNY8Yy9dJriXN9zwqontPMsnOE23MIYubOoPbJdSypCPOT
XKaS2a11NZ7D/osvy2OGtqFu/ZZO4VA/RKY3tyDhMvdKmPWXzo5Mk04tZHfFF5E0
74AwzTpK40LRAb9bYY7a691wQ7L67SR8MhBuV6Hzr2MpaMzIiUWXd6s2F5kyXX+J
flrAzVaBCyHSeIrLviDEvL3S5noLgHhYo9OjFHCWJmtPgcWMuJlgKWQe61iuz9+d
tE076vZXpavqGNeeqBymuNmoyVZEfjKTi63ShrC/Q7Ak3bxPzIJhU6gnJLgwPK3B
4izxskMMSP7IhKPNr0xdjdHdwutBSZx6HrnbI+/Es5swBknIrH0p+DBo8JKS74Bh
A/HSuO4PhFAZFLsW44tOBMxbDDSKlaZx4t88jbDisEbfhYRVtBMgUzFDl0DEXRBY
7X1YS0avz0B+hfTapMX3J31+8zNBmRxH1k18AETeYE2m5/ivCnyvdlAnj+kpojyK
NfWJhTLxrqhItmb6DQqb1uFzYgvcKedKQj2R9I6vqWorInHUffjOPMS9qBqTnMdB
hhiFej0KKQlVZWCU1X4uQSpdP0Nciz5FhjPxRaN0aDIze4rpZVRGr+9Ss64H4XHA
BHuA82UQLnfcX4bhyuQTffFnV2wiiHQ3TBGrzhVpdFrvNCLd+fLOQmRpfzZz9C6z
wXvMM8xH0XKe5sszVOFfw8DOHI/WxCw4fT9rjnVQgw8rRuy3cZrfsG1JCJqcPYsZ
/UyPaoYm1rsmbRdEMrkMMWFFbFSudCllAkWjL6lqkn3tDKGXriS8DfODt8HrYwZE
MDeOSPJIVJrNmeFQyEqkTIgs+pyeBz5Y7CN0yyIHXJlQI/yk6aUmtvj/Kx3NAxse
agndhiPncOLWcg3lhSGaXYzsP1qGe4K+O5Td0zc6A6YcIjnzB1GOXvRWbL/Hj48T
GdfqdYms3fjjlZFUPjHPuePSznX1EZpSfQCqhxr8HUu+YHr87MmO6T/x5QFgnXwt
nY2+H7pXrlPrxqgIJptFwqQWzjzbB0A1fzpSyoy9izWevDQImCNgA0T9jnTvOJI5
zgw93k9BJMIDX1U6pVopmKgWt6drXJlrGRAC54b8jA1VrMyn1I+f/1OobLQpm+ZD
WGPDkqIR66svfIhiH4idYCg+fu1U0oIElWqLAnbZlkCrESngoztLIv4hW+U5ObDD
HQ6wzEWJSqgQwkMWC6oEusLVIv2FNckiymC++nvE8by/pbUOviEYGxjkRrXM3k72
h53Xw76Lymy3U5c7A+D92EtRyZPcOgFcMQzP7WudiaWcDWrIOFXcZ0udc2rQ/lHS
tokG/CpVvVy83pRvY2DgsudLhlHc1trpiQscowT8cl7ae2eAXlHistyf0U+Ju/Ey
oOcPbDE6l5OoJS7dlqyYciPUHONNv7MAOpv7qsbk5WK4zWpGMCgDUcHjHn2r9Xyc
biooqhwfa0w7RWDQYgt571yNSrzVtEh6SS5xri6QuqTlD4TvFHpR9xvas5Y2jNfw
9AGP4ang+36kd2Bs5M4dqiWEFPkdqH/XyYOigHm+50I7K4pCfkNevtiebPesewiZ
yyN+DOZCSoLbdHwAuE7V8u3Nh5zjAK4FYDUhGvMHFf6HR19p7aFaLXSZ1z9483XW
EZaad71FFhTP9Oj4NSzne1gaMWKGbhwL/0N1vAD0KuTnAVtUldO44vx7aUpwXijy
aJAfd0PLY1+oKIz/Ig9rtmStQVfkX7FhG2tSNeEoSHGjcrCnrSAS5BDbjvCjhrjj
izBRpBg9mdoeks5gU328Yqiud4recqVEDAkvStyNvEg9NenmpnBy3vQbFfCJ49zC
DL98C/lfZP5YngIobs4y4O201pZSkicJ2MlvS0H59ljDY7WhyoSoioEqU9+M94E6
x/QiQq/YpvqPLA/WCmRLC/sDroT+/Bk329Sg4PKbfON6YuL8NkNgF2q0DlrPbTA9
79ARR7N9Dk6RhKHpT8zwJ2fc986crZSYtwh/r/usfJf+wyQ0G35r1X+r1P8lCt7D
IZdi8W+OMsOXSl9iSilGYz5URq0s03CEwBkTTRmZ55lbguCNVn6DSKWwj7PlLGy8
Lkuj6Mj67F+4b1wco77gq8bmdHB2R1Ax2/w0rNR30llItcJR3ja2TdWKzAA9wdiY
jgI8OXbj3Lt96c77Q7G1Pox0uC59WwbVnL9rogJ5+q0/0VE2ocJnrJNOIMrv631H
XanVSqeD1MQH1NierhRw6Q8XiOzrvS31fZsOqgMN8sf+488B8HyljgUGLnFy8X6i
hJfEwj9gMkUN8ZG0eKHuaGliQS/fk6Z+I65DUj6GzbetcDFK3egBrpcf9WuhXAys
+9eNNySgSffUruiEP5PzdhZoFc6G20rJNzMvlMhMkI/tQdPZMcrJ4UzKwjE/AvsN
Hv4dMLrQvvTibXeM3rJwwJQIrN+1/rA/S9r7IbiXSEvkPKuqy+DS5Him6Yt4sXTN
4DmJPonzMy28cdmVe5yRoSgcnls+kPnAwqWloA9f0kFhvdHBtwE4GRQml8US72Tq
nvfPB1Yt7szgH/NFpJFa9l60gqXkmIx369oYaREzWfWiTmGV+P8JC7LrgUL3iaoS
1qp+328hXWiC//2JGcGw55iQPut2dOQ27Dzto5p10/LQcnQbdTUeZSOHFhOAdMeb
oPuw1p6X2Lv9uNkuRZreRL543I28th1h7od0oG+8TLPpcf5ylsgSQu9dbqIhaWXJ
VSt8TusIc4nAQ+0Kp9tyarx2fr9PeIh3kqKRRsGgwnDh10QXbpF3f7um7lLw+h3H
uJh2uSumMfexA4CqSmxG4uFTX9pQnS4R/W5toGBQeDQoLzxLwTRCMtTVuJG87D0W
4s/FK94eoH3hyGQU8CtORA28dlhUMhy6KIlfzL7jgbRF18tv1yu4nHevLoH8Bnd3
zGVBxlsQCNYbBnC09PtQHBGZPMfw+22hIeS+vGscPgagPFz36PjJv5Gs0SxpDYn2
TyTm/fbaVfQVzItO1msfpgvcBza0aVpg7mBKGtDzIu7CUsaW0jGB6TPcjtNzhyT1
KXIeOQmLQ5AaGNRnRt8LyDRflRKjTB3+OU6cxHdizy++oLQPQNjyqtGCIrlxlz93
b+sv6vQRkqepvDo1iW+JzRljwiFg2LkrmIFbnPjdcE/WAGyW8GEBvADVUrCl6pvT
20gZPb0sFHv7QZIQh0IJTzRVuNa3r9r+UWthAaQPfITE+5fPkTFfWAwvBQB+O1Y+
8FxiScchugmInz7HjYSs2BTrMCmzgCN14+cCoZ9RNitGuUAq4kFwiBmeSs/UQoqJ
hw8/IXn0KD4x0eUIUjDqiKhKu+QRab3rrraPsUFVMB8xbNZe5o1ijxbyW2DNRkWv
KBYqdLBWXKjA5XxRA/6ExXVLCnv+yu0QZzai//n9ula47aJfhkIgKyYAiYNyB3B9
i9EgOKgJtsnrCUhF2QgiewuB5IeYhECMIbBisi8eVf0A5r9JZO/W7X+ocu1S6l2y
zAR/Xhyg9CKEIljjhxKj599jDBeB4sXWgc3ukGWR/tIZnYEHkynckp9ijsaUOtpg
u2wqiGhneMZpW6rx2FTTK/LerG5imnoJBKDh8RB2/ZNO3Qb4LmSrhaMfteXS8vhj
aQRWx4Y+YBwH1NOT8jQPQqX6vjkwrnzgpddHk52yUGUXsohJ3glYGIOkoLfnNzK2
QVxQih1d185W611W9ZnDAa70hx6q5iM7Ewn4lUb5Mms0XrOv2BHnIxbOW9sfCfhc
OrwlSirmjUfLmq0tqwSKt1/hBEHgEzTIGc4HkOWFdfe+W25g0Fk6lcfMnmHiOZdg
VVGaU0Mx/yhrJIaBpgWOlUQXmS0P8E6/PC3dNKXT4AulYrBQ6nwhewT9MO29BMp8
NL9Pks72aDZhfuMERRz0XqCwPBIgb9KPErGAn7PLQKkWALzMTVVfeFDN/0f2zhCN
3tM0RM2Q4vhZDlNz3KlikU8PUpIO0zuJ5YdmpHGnb1oSXBD+7ZEkOjpBvka8NZzV
1P6uzJS6GIYyGTx+rxok8pOEg/CtCWKXYW8HFPw9X3Eua/5aWNM+1L6Q9woYN60d
jZufryK4cXSMmzOA8OsGuxJsEA/L/8B5kLj1erxNWcKKY5YSum6fn4if2Ravn6QH
U2igqxlYZkY0lTG3DjbfV0ovADkhTgABoFQk8SUSMuQt7WFPZtYx7j6A44LOCBiu
yvohKUCUR1W8HZOzdJEhKMRsgEeUWi1OJ/oXoRSTkaAg2qkxahnYV6vuX/QQhAes
0SGPduXD10Wl1cXMaq25s4GkBqpAaqoWQUHeBv/pze8cx024An1pzjXVGKj6A9vu
T75OpXOE8MD5tCQaCkkIV6bsaQ46LzJcvzgd++XreV2fmCFuwu4TjDqzAVVSnOFW
8K/Ddd1UkwDP+hptQxrrzw/j25sR3Kv8wdD8LEbn4Mi9451WZOsCe/WLWGsMZOBN
ekdbzUbTNSG7ewTM/erPJOcZlUK40b+Rvsrwz92lJZeiwNRsTVvGykDo9kf+2k5u
qkYZmDVlatDs0ZZ7zsA0uXYJvv7MpbUOSfSOM2YjPC23y7+HK8tgo6mUGBQFPAPv
+RrmNW6K4V913Wa5MQIeBSDHNpgZK6VMwzwkgJ8IEM8MJgqr23/AiIRt4BFNJrO1
Lf9GiPF45O1x+RJmN8+ZX6bfqlOBdT5oUc2Nkgxwx4RpZXnTZvgWT0PsKVRXqdMw
acrImYPjgOtSXCsl4TqdUZ8M5StfvGNazc1M4PI3Bz96FE+6qTPJJZ1KTB2vbBoU
iNpaCoqwu/sprT3FfBBWZ9PXeB7ZmLAScPlAkXAFZ3LMht6x6cyAYfjuaj049LIA
nlc2L4XQcjpqmrRwnvYZFNaHoUTtC2NmBz1g+SI1qEeMEdXeHzthnwip0vnXRhNs
zvlzeHB2ySpAuf08/Bg0hUUIz4ZJRe6ntKLtpI468s08Ayt7iy/8xiSbrFAdgeon
U9q2SHi+pSb0C8aNFMkBs8ZliKUWc7KMJw0wmG7s4i81rsu7QhFfDb3G68HhFoyt
a27TPvGhlDl1zdzBnbFEyA5INrYhoRcrpl8ZoJbjqqtOqvHvtdRpYexpJkoSic4H
rwjGdWUn9rdyHIyK+WkuexWgf6tPkumZ+dgGhnyCwDNvyG+ismMiOyMiU1fpmjc2
8810Rca8TO80cCLjWfHyJ5ImY4JS3V2wBz7E0HHIs79dO+GAyco/WUbxZryQJ8cw
hO6Cw20CRmWgs/nWhsDmbCBo2nQPBoNyHjutdJ6z+w9osHz+A+9o14eTDQshocqU
OSjcf8j7goK2T3NwW9vybbkJFM/Om3lYCchJIeEtEJqCP+9nhpK+8b/W7qDQBMIm
VE2DO5KX/NCI6NCn5VwhSIl6wplesihEsL4rcDmbbDkbrDWIAMmIYVeGJCSOVQig
J0gMpA8hON89UVENNo7q6C0bnzPDxkDdooOrU8/Wina4gkud1xrXCfp/Z87MKWOf
3PlQ2hxbnRKgMJn+SlV/Mr/1oEJdy5Z+shKU3LpT9MM7Xf3MhTbm1iR/tPOADgIZ
`protect end_protected