`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1712 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
4PLO5jSby01Gvgd+5+tHBMMkzXSdNlDCHPVmXX6Wmd+1RiQkqd12yMfPk8z4cNpG
if9q7MwEYndkbnYVCC8spxblFpKsll5DYC7nquBZS2ldfIIzahpjC8fE4DKuIFqF
vdUVAb5xOt6gk+OoQ5e+LL5Y4eDs7O1x+GWG67wEc/FWpcxO/LknVB3Nb+91W06I
6ohpFlPJ3Mqe44ZFJyGZaZ2vxX085ucWkTwp0EvwLDIR30xlwemMZgJHzluHYZx1
xjMCl/NXEPPigZ9e7q922q+Cl/mslQx9DjyOXg2rc8lsLgyIzOiXy7q/NNnj7hbu
dqDl4kcDlYwtdvzQEvTO0LoAhkhiIeVCMNiE8bCopP0Vp+OdqRNjl92EUz2yoo9F
tw19tWgBvbG7YV5zAUd56iMe8vJdRg61CWBDa4U385pNyJEU9csrsDNjvr84YsSV
kF9ajCffhzfHtlYMRIakDRgiYkpbI2rRMBGVMiYL9fKPSUrfqSkB/BJu3aY5JG/b
rpkqgwMomWGp0i/RqXjG0O30ZHS/IahQa6keT5swABzG088LsZs/gZvl14dLnDrn
N0N/7wIatc78I28tbsQjlEnnaOEaq9BA+5T8sCm6vH0noBuBBPf5uvi3nAHoNR71
J5qyf4xJCzA77enaIdDU97SJwFfDX3mYZqi6dOvzglXoHc/OBunPcVBnT01/Yy9e
edaYttaOT+cGLrUe1X6+ELQbT4WNxFPmItcrXM5hPfxBKtG+nnDj1SP5wVY8IS2Y
IflTSncwOwTk+lFHk8czoU6r9WLxnHbFhd2oN22/Rqe6X9FkfjtYSYZbIQtY+nuM
YzI/3xf61VYq843CRX+9Ch93A12BT3sSjDCthzzf8OhDxGFWR9GdAeXs+12B9ZaK
uGSljgv65Ggeke9dhGWDdTyWOWZELda0N5dPPltbspR6OIE3DTbbl38xgseSsMah
6NAkrUF/QYZczooKSZyBSqAvW1ZEbT+piYlhymyE/muBC5uD8aLbSHQ0gcBFH2rj
2xz+EoLL3TwXRyWCv38ZUNMZbBYoTGYaK6uBOtS9yewu4H6xKXu8cbx/AT/wR5Dj
rRDqT8cprLpU7se5xc6pod991TZ2meTy/M9L4Sql+hQftSczDYVHesRtI1Yf5UIA
50F2XPlTmlRuAcQ/PTFVUNCTZ/TqlUguXyAEZ/rvNayBjfnQAMqkmpyM7bTUkwKN
BzJdWA2Ns07W9sZOm7+EzypAeKGssTGjOdECmtRYpO7I+CwVDPzMwdiacAcj8dnf
zEcPyHowsPbqdBtTq7oJO4nSiT7GCe0mfe+X9Z95qHCL5I3JEVjUY/fR6dSEXVWY
CApTeb2UG4RmrgiNswEuGrccyh3QECp4zxv03iE7fMT0RuSTPJ1XslXZKEI5dvvs
PPFEIoILOG6xanFPKwTTppaKBGFKnJn5CkhnWgezlRrVewHDh4Q0+GaPVh4SiZIt
1oaKAm5N4GSQlEvRRGyBj5pPnX/QEfnIarAj+c4pYnYn0LOP4BOQWWuN+j/2t5z1
Ik3F/l/yY+he2APfB1hzATcU63EvUozB8rnM6lWt2FwKaTvoxn/uzGLw5R/04nqr
Ph2sRGIC1JCIezW6k5Cs+OXVyAerGucEBlLmBfD2sHTeDUS5/Zg6Z+dfD0zBVLs1
D2yf1bBphSDwYUhDH+wuaeo2dLFNAOxRFLVKu1dcTjsEhRPG21zSMSTs8KVMmhTv
yizunT4Cfr6NmtVlsOiXWuPhyTZHa94umqoYgeHHGKR8Ygu8n5owKu88FyyvW3z8
HCFdTJsaGqofE6YWmJzgssCVdHPNmpMsQIfgOnzklP836JnM94jBMxoX8hgCxOsg
A/inHPuIUE9dnWKI6LcAF+mPVf3eOpYnKUjvcSKqU0jYFYaQl4F5PPYpN829VaFy
DkLukCZKxpSCW7tJEs+Z4Z666G+qTCBywjgqc77Bpd0CmjaIM5i2EPCrZCHBK6HQ
qt7+pJcRN4OtE93ARjEOkRyFNgDOUC9ws/ABVs6CgAiJqdsXafaICvWeHs6Md59H
GohhjqqaQHK9rM7cxIdoDiw5UQbVSLIRtaeyQnegv2C2C3dBY86dbOp2Mv7NqcT4
dVSV/h5eTRjoNuDoCfLy4WX+ExH35s4dt8od+XNAfpY=
`protect end_protected