`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 34752 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
3JbtNiAekMoRUw6FSbjvdFz2Eg2XxDLqAd0CkqhFD4uNZfdtVY1iS/4GU9ADS9Rs
pDdnIS/DUroMRKrbZ24maA40kIqGKij0Lr1kkOiztB4VElibkeM/haiv8mj+smMJ
1/fpkFE8aFSGwczxCN4LBubHpoNE77SfSRuRzGXx3U5o+G8Dl67EwmESUyeCRByi
8uxFN4NfpnqrQjYvaOCsJSR08470eD7ZgW8kY58+b5VOXwE982LqfxxfnO6V/E9L
oSqjdHxPhGLSNJmM9UYWDp60NnIYFTW+bNmOAhqPnQtqWv4hwuhN4wYr3ngfneGN
xWjP8/MzQrj0fA94UBkjiB6RhhA5Jbt+Hvis98y3t/Wef+BaYWWmCnpKq8pH8ZuH
b/ad9nMGe3bwcIerV/oc8Ew+X0h9UWr3RuxcZ2mHTH/59rGuE9JWMfp9Rg9Qk3tM
k+FPd5jOHDGjbjA9841NIQmAAB5KbVcCugG2hsgDaEPxvgenbTitQJFvxKN+rUTm
IX3McrCkVL30Ng0Wvu0lEFzi83md4sUGz6IOhSftuxvM6YleA3PpqGRy3iSJqjA/
AtJCk4tAfdMdSMSu0DIOCIsKy/GiPCC0h7gF1HCGvns8vmQtR0Si/dPJnoVsKqw0
odw60d4eqXvM5XObz7N3QMJemLWblmSnoBopYjv5flzO8t3go7bhxlxvIGybNzQk
X13ZuGP2z8WgSallZUpn3BIjjlVOo1djguQf8/YmgJLqcrD73mXIc/IjF3IRuPve
RjJNDswG4eX6gVgT8Blv0hzSrHPzexwO/gNr//j4ekNsMiFBrXvp4IxxL7N/SdGD
KvMPVJ05kKIgCNMYrPP3cM7dHLKcyNE9M5hgik0xA5aYUuAFbqhCfkQUSMRAXe6j
ymA/BoAd4HXu5E9PEQQfeoFcLML0XhmnLh4L930n2mRZ5NQ3UtfZh0q/3h9016el
oIkO90Si1scZNLkLPqbfKou2gJeuuI2iBmcfui/p6F5G0ILv4dg+1bnPJ/lEjcOo
ZAGGEPSUzmOh1EfzJYvJkPdyhb15LUMLcRanLWMk1/2h1WDLvy+Tlt/I4w7gOfGl
W8Oq5Lx3LMBj60SZGyxeHKaQCzOr0GLDbmU5RJF1qPyUZikskZdy7dkdn+zS1s7P
jXR/g45vLtHab/uZGT8i2PcjgBBKQLe8cIyETacm8nB9BysSrREJCxKdz2iXgApq
8i0JYdWuKEU23aIeyZ/a/yv0XrDVPHwdWwK5teXWTgTL045bdh/4VHUymwG963Ak
YPpx/RhaPV5MPAt96clwiiLuE6gTg+6nrLDVNW0kZGOI4U0hvkoaw5VYynpoPoW0
A1A9F/gVYbozwxOnK5N+mpU0sJEH4OFHwfWcK12Gv6xzT44pCj1oLCORAZdFnsmF
z39XKvccXuuqYIlEnrpVMYQRiSdgrp+FHHn/FwV9GcXOhAe5MdNjMYbFkoma5CKV
Vx1UC7PYuSOjgtDAg3IYCd+gb4NRBVagOfysRh1EqCWCyaHsFR2XhkUddxc74gnw
9fuN8giJMMdZamxgRMI3+MALpd5yWzS6dYu+U7tbzQNYOy90VAuWhvGdlNFRjKQt
rPWuveActU+kZ2LIe5CtW7cWjRxVAaOR6NE8uQMledwgH2zTaer6sQAhzrdlgCZA
TGjqGzmpcTMCbThR/1GYunOsuMGTzDx9oSKgMYzsiAOQ11aeqjXiGijcYx+SD2nv
3xJJHon6WFkjETazFoK12NULOO3OOWTVELQtNlBURP7EFEK4XG0d3z0oqLdb0Pxu
26Qh2gnYvyTZsfLRbJi2zHoDAfNw2pT6W2dCXm+gMHTtaBYQl38G4QosEOJTG+PE
/x5bbm/i9YGaWkbX/Qo1mYpzoIF+Co/UjyKz90IgptXHMh+h16WYi/rYGD49ac1q
0TWXc2NmwDm+2xjRa0EGmGo0TRF8DxyVOUxYcRvRi7KHP2N8dw3osCPktZ+FAEHI
JlgYRUDShHo1pVeGHsjzKaIkKoSecomKhjtg9tSwhfMEEnilA6VU7tWuiKrzx2xk
/EDzoiYcac7m5xi6azxjoLTYp4OqqMy28lyLK/4V04QfPXtoGLqL3vao/c9eerd3
CVwa6dpq8JlDCcueJPrA2n2u8vWah+wlUBEVnFqlZMnY4LIaWPe7AjD0YZKDv4go
bwLt51S0f2VMK7s2aE12lqZc3w7dSN9vxIDjG6Hl70ewPN7krYBpl08M/LeNcbB1
chpkfqOOgr571u1YWGgX+mJLbX8Lh13ffqObwn1/Sns5c7gACWfHqt53Fp1zS4b0
qfS9mq971vcw2/nrGgVWNc3xiU65gEIGyYLuTRthfLfZmlRN10JHVPDE5BJp6byF
fzc4XzAnKIMyxMpFamwcl6viVDcG8cbtYYUj0TSW4hcqSDVax1SpS6gD6mJXhMXu
ZlNrIPiT89xRkTwT7rkfVhZC5mBLBESWpoyempQljYdtWl0zyfvTWx0SzbTBS2x0
NwSnUKYCdV6ExTti5zmT2x2BoFQtXum3dY4lVXMiIv7S8xWP/vC+Fg/bVAPnJvSY
AFX2m3UfRegDeKsJ5LIapZsU1Pj5CXpqnOzFBd7gkM3DxXmflu6V4zdNh4+yR5uj
O7JCnPf7x5ThIR0OsDy5gU9FTglb/V14OLSMpYpweWyQcv0Q3OWb8Qpo0Bch4S6U
pxnl1Io9je1/l8YChfp/DWnzq3X4YpRzI97f2j9VUBmOo2YT8w2quWSRgpvip/Nx
KydzDnb0jbBHyXa1ijBcps/5qc02VqFfrhK9aOgi+bTWv5j9hDo412B/Z2PGhr1Y
4fqR4ecD9vKgJFHQPLsoIjO9zktVw/vP5IAvE/SfMEkSnUY10an7suxm8zdkIDv8
QKhnUhqyVTdP7D+tr71xdi0V2i4W5XYjBk7FiTLopUAQIIIR5s1mY2H9Bs8FGTkG
DH5z4L7Ai4g4XbVEeVA/xOzu8YyzEMScSx8+hr3mLnuZsPGlqPOF4leMv+q4N3NU
HRljHKocKfqPdUt1E1oBoBsMJ2B3/Nj5GI6b2hDauj4oG5olyrFg2DI97NL6sN2b
/K47mysNMgWzrFwRY9LvXTKqYEF+G370NZrB8elJaShL50DrraZYNeDGJyk4MkbK
BSxIaIqdYDjf/fYVYiBmLVIdj4lcjr8gfwE5gneiAhTjut+pfW/7CNCQPSB+1z+d
4jUYIiuEAnmeHtBYVaIv5hm7CC0LO8DgYLker3v+WkkfHSmyS8WDopTCIFdQvbi+
O633yMSkYIlxP8yTawztLDnYEH6JobqfAqyNEiBRh1Io906K4Ecd4kZhCIrao/9j
KiaiEFdDhZsds7aTqW8vC68Y6lRBD1NfbAcw3u49wP8NcZ/KAY3w9Iv6NYmqkCe/
QYARP1wYk5vQH5T+8hfVD/YdQmVXnI0D7/9XJjZYyexImBAcc8p81x3d3coWfovv
EOJOtrIQjVvkYtbrE0syY/o+uGFVmbFh6MrAyzRwK/rDvSsLBbIW+D5BRq4eYQkw
hp7UWJHGJp4fsBJbMb/CiaSVKqLPEdFsqvGAI/npMYlpQD6jjcigQyBPVn+RkVuX
qx2kfOYiUhtnv/pXFiIeGbLeFZIaq6V4fgVML62Si6gSWjw7rxRftTZDqVgOffuZ
G8cfXXLhwt9fHXnmmBli7ovZHkQ/y32n2waTQQNvcfptVONs69OcrmL8Gq7rH4ON
aw6YN73J5AIiH9g3Rtc7b4nCyU/JCVDX+WHpuF9xWXBPWPIEN0kowDa32juN06sH
CrqAKi5+E2qCoa76iZzSPMnpZpdu3jpDQ6XOPMBjFacZS2ndLxXd6b8utyAh9RFb
3IkzOtQDYGzWSOIuUjaCJHXbxS04YO3PKC7PbsjRjGxuPLVPo0y5j5JLAHl+RFyQ
fk8pyt5S55R1RhT1huKJnSU9y0LtT7HB2QiZLN2V/z63gY2vNmK5EJqMFkBzclor
R59uoCLxKxhl11uAkefBw0/RVR/3uTF0BP3mQ79TDXWJ+RuTys79HPNcE2WD+Qgy
+Uq3z4v6FQwLZ2JOVLC8BXvfTyosdF4ATuiOMtk4lJO7k+E49FQ4IgpjR9WfGl1r
8nufIXtajhcCynyR+ONdDA+4LeMX1KttOK62S8GNh9YI3l32a34e8B8iOF9nmR8l
evBIhNUDtow69tDZyQkVdY+hyeL1wsRh+ki80TiyftoT/SMWuvdcFIGfJixyVdQc
L1ws1tQzTY53z2ROCOXvrY8Om6Icyp5pStSSTf2TjMvFHvMT8H9yj6D+KB1qmTwQ
j9rHsUo8otCbmDeb/VWNW9J/QO51GaAVHuT5+YSPlFdRofYxmtDNmuMWF7+JUBxb
7TO5mfHiHq4X+M0UhoIgPr3/2kJGFbzak3K947ulAZiXl0rUPgoG2dxzSc5pwkqW
NPh2uuCjKIBxayzhOHyNh/5uvXuF7AWHM9Oo3U5tJEIhg2tn5/QqT+IUbdxeowF8
Q1+4iQqde3aQ3vfzu3Io87cUmfbKLBUUj0y5rX7Uq3YnG0DvzJ9t95rLD595Nncg
yzHYpLTRoLXLN9radTNZtgGONgBjnUbeejNUbAm+nTQX4lO80sbMc0xkN9XPc62P
eTg0fMCyBcR6elwyCZEN9x9tBmF4gwp73MKifpWH7uhN7EXGWzNYY1Osj/GzGCyE
sb7NBN2zYspXmW6iXpaSo/ylMBntUdU04aKMBZ/ZqndfQnpLzHxHfDbjklD9pev+
pd4GVvWMj78MlNqEIO5EUxUIKrAi2K32LgXpxnLuysbNr09s9/y0oHK/UsGbN8MV
m+6UFLm/6ytwlT9Pew5YGbWoNmZ2z775l+u5Ly5Nj5P9CF9U9JVFnD5eRlGwkGP2
OX4VSB0QLLl55kFHvZXG8a3sTChmLdcgrTTFJcmKlAUK7UMsAelNT+7ZHKaB8UJz
G38Mot3q0HVrcB0s1dyz1SnusLPKmwpnlbLMLqy/R5X/cMs0bK22g6HTI/IBrXf3
6Iv/BlGidaj+a7WPD2SdwoWLg6ucP5FMSTBkayrVYoeUtAj9ZevLbskzDaZib7Oc
bRzCallbaEdc+RuN/MLJO5GaLASdu6/zyo2gcMYLYMoE2cN7kTV6ucEJDaVj9HD3
s2IifhB72n0ZQ8Sa1AHiFdMuQOZ6o6FZdMX/afGRcC8Kicu/vfdqlRzlvtROzTWy
vXThQuTV0tpSf5U1tfVOJ/dpi/jDCiJyisLWzhYW/qIRTnHDZJVw8MiLDrRdPCkK
McwMOe9vpfTiKI9MPwFHF59CR8zCYrIzG3Go/WsPNbmEjZYAiFmLqz+Ry2nRjNrx
TET8fuK+BWYRmGlz3sArXFcDWKhoFSYjngZ6ttJtjM1nPiHfN2CyiIUi7arBnN4w
pXjhNBgZJ/bu0ktp750DLDIZBgqQNifSVk6pZFiy4rNrDEmeCdPYZ3Xl7joPHaB9
ianF+EMOVyDSM93RPsWITqvKLW+f8q4/En+KB3yvVwiuIAFTjVTPbOaj5SbLUFrG
dnb/LpV2OizienRHVqJ4FF+ZBTBpPqd6SNKWgszWh/T2/esoL1zZTpUgbTU2YQzF
8SSHtrvYeuSvzpsHqUg4nISzzNoxB/iwGv1YXidAeW8UgYDVlgC9U2JAserAzhm+
YAYsY/0jfQm8pgrXaYRaW5z5qaOtOUE+45KxwsBjYXZguv/wKz3pumb3wqbi/MfC
LGU9NsC3LEQaB0AOtnLvWr0aIbaDk68yeNwbEQywieglMtrtthPO00Xayaxp90wy
ISVbt1ziRS3nUUPkZSnMK+cbmwgD8Q0bYLBvwWxeVRfjJ2tmrMYlgDxOPSfI0s/u
bK3rcju1sRzvDrlaE5nUkCqU/wuaGDrkyppx6HUscWZxNhiXnU+9940l7F1c0+rk
I9AvqocA5fYmr48OdhSCNEJ7fY40m9psu0QJeJxnRbN1Xl9i4TCaTw+Y/OQXdUiX
99awgErjv55BjAINpe14Z/G1dvzFvkvBV/2B8E9GDJc6BUtBsefYvcFigiMEyVM2
2ADHh6goXuVwFdikFxSy2R5sbODizGKBoZkaOzvD0zQQawHd9lztgZzD84KWYYE/
nCrTtVz7Fz944RNfXtvzE5KnShpdWNsAwgjO+XdADi/tjy7TpQ7cI1nPlaaZXjwp
Xy2sGAtWSS+ZQ9dickj+rdj3oW5QydhfoP39AdnZWvHORoNoWHdhx4y3agFYOHuH
HA7epdl3x5sNLsOPtUzt5ZancqG/IyD9AkfTcQNouyWdVU8r2mdXnaGI6GPLD2n/
mpeCmAb1UAj1rVoALPeqG7YwJ5SHCb0krivnNJmQY5J2tqaVEdAP3elVCw2D4+E5
S5u7e60Wsz7aEKF6Ido9T5Rabeid31UKtfrIq8ZGYne2xiG1X2n6Fn1grhKxf7Uw
k3D+iK9GmJKm2eAsxzE5dYnJtoKq3tD5dN137TOvpgTB/NwdiQIkgvQzHkqNm3t5
1OD/GZ+cD4IoUdENLa4FvmRmJcvORvHNh1WmNko95q+iq8ATK54FtQss7BplMiQ0
eAS4GQKKnpwQNfecLsSGRX1GMQe7IBMguHZ+PjqNU8xfxyNqfwgK3tRKqvUboGgx
8KvP9fEY0id+KXC2H6DyByJSD8eR3Endj0CveU3y/M5XBItkJynxRYpdm9LbuEsC
H87H7kOHgs62WVs09HnohmlUbm0U2WBRUg3kdYoRe2hrVkLJybrgbQa0zFqmePck
usuClXNFvL0L0vmNLzKr08+0wlX5xerTugfBth6n1y4HR9FslFAUuus/v9zzE4od
QB57tJEgIw2Ff0UrxsKSEWAyjxMnPvRvmbp6yHqQze//hCm0yyMV6zjc0SlqE4Ax
VQsIs3JNC/reGcnadUgiBqYpCM1Hdb2kbHgH00ZSdqINtt9JaEEPRgJJnTGMoo8W
Lyh+dxJdqbY5oHxSVdFzZGEJTgIm1CGRkUaKuXusWwlPLMdmGEMj5Q4yK7bJf2qx
cSPoNO1EEUNendiL0ragSTHFexYn/Q+AeV96rcQi++ZYAP7tVMcIr1tRpOOOHPUW
X0TQFEVJ2DHrqIi89pUwcmbXxLD3eeBYLLmU3KQTNRt66Fd8hA92cFP8VXsdsa1S
n6p4X5ICqYvUORUzHMHc0g2uis5eQCl4TD7k44Byauz6tyW7wBvKIdetlbCru/2h
bmWDS4XTSZHzuZy5il6Fj+rnXqnwQKSI5R0MxHuwPqGIZDQhv8G+wpTCowwd3Tx6
Mt3HtCF6rPPuw86KKt3iZkpAf8Ib2PplIgHlXsFc6IqIm7+o+yQGWZHCJgqjpo3O
PQ98SRddmG85u7XAjw3xIOVS5OxE9fvEBrFlQCRru9TcTaHhA6/JNduXNBkmMAuQ
HxkeM3PDd6gk68W+FDocmgvG/0JxcU35/YTIjiR7NBHZNP6wQ0AofD8N3YCP6XZY
dchrRmQItVOhA0Hg/+qK4jjeF/ZVc2377IH0/ORWPkXYLjqxFkonsCm3RUHOgz9n
zW2SstQjDuzFDld7/cQ76B1uAKiE6i7FsAy89zC4nMZ8yPksDOsBb5nEt7hOGqlN
KY8UxIuIob5+fKX4HphXfa3jtF6r+K6ZWs+vFLhuRSf8WpmgYkAMOeKHqbVV6EQ1
P3NYXAOqh7jJrwWdHRP2kC+2Csa2F1iyye2+fTvXwN0AVpjKUNyALn/BQRZQnvKp
R740qGeLxf0T+vy2v0si+/3QXVuxoYCEhsa39QLok/K4Ab9bI0aV8JRKEz5cgv91
3fpTw1C/aO8fCY9/3eGzHgGP+yvGv0/iVoaWqCrDbG/b2QqiVcRT3nglSGjnjRYk
0sYMRYPbhd1oe9cJ9iMnNWaljfGFrq9PzN6dooNsoc5WGua9VmBS/uRfvWd1Q7ju
MqWCfi7i7YpjUYEFNIL/Re9cw9zWdtw3WchnvYcWr2jLeSP0rZaWYvct831+VwqX
a4ciFUmlAgAZgUgBOMwy4BnQBh5TPQJTxDMbPQnTx5rRy70WU8/p2pY/ql/YFm3S
sfrCAgmGDMA64qIalJYXClHkg1g4igo5pvRaSSmUApMwjSLRunnobwQjzHA1fhNI
rHqgPw9sVyuLR5LYqH4EXKBBgh2IaZs5XROoU08qfPqLub+ng+Irk78//MZRqxiQ
2O0y/2yPU3uJJ7zvZrXPb8kWR2LHWKEPYSl+47/Wk+FPf4J0Y94Ayi+0NiJuZWEF
PzP8/scMjyq5a/rKNXRB93c+mHGPlqYdTXlz3+2Be+uC/djQ+eu769VU6aOiYttV
ywhCW6tMVvyW9B47eDzq7+nwrcCDuudSuODMKmani6Ca+MxGmB7rnuOEnP3kWxSn
OO3F1nq9OB8aj8JMhxJ7KNgRzbmO6IYW8MIFzj0mbOTkHPasGcP1j0ocAP71w4bV
NQdTYL/cog4vTPmlAZxq31HmB9e+pOcCYXcF+zWrvulNDXacsUvQdMBIF/BAiWq8
LGfLXa8gKOTzemvGwIukuO18CMfObWQI66WRgZ9oHgUsFKi2eV2cXedJhO8CczyR
ynTYkAs1Hqry1jODudgKXBHEPi4AKVHWadg+pMmXibyCodY4KMTut6kq3vNzj8fD
tYtgIWABMACHQbQZKyx9TqVCvcReaxyuy5eVTupcSa9C9WUd6SHtrLCQOO/V/RDs
OMMyuls1F2Gjf9WMr9/Y2nAB2JT0FwqJfnVwDsmTuLLNPJwaqKXYIX3GUegrWrzr
HRQBwU+HL3ZPvFpUhXPEqvnRTf+zdeElyfUJhGymbC4ealnyeGF0slFUGgVMigik
Ek1Tug8JWAUgSpTjfs+aw9v34GqjI7tYGvd3qfQ1iV3o8+CyUnN7ZJUDz83cGv7N
m0+hPSfXRclyi47Lg6GvjDyblqJxANO+qV2sYW1CJW9wzykjWhh9gCFGd/64ULAm
BSH6+xWg0N8LOdwzHY/8DOS+tjpj4mJH6ApB3SVqnbj4XhRmnQepYd65DsFC6Tm+
RQxVdn2KTtaBuOy0JX8c145JXqdQane7em1GaYgG8AMFcYuSRymZXmhHlCW++eDb
9vDct76dkR1nwgpUT8dVZwVNTJ7hv9Nmacs+WOb5y8bFqO0xa+elFHRFmKswG12e
Mu8CgpgwNZg0qElPQ3j8XzXIlsZyPCJnTYotncP80fmGeiMYfUEbtPjCKAg384GX
BUR9/J4HlZjhLKiLER3EMEoOk1F+6TuYyFYzrH2PaRwuOUhI4+KcjnDW1Ztm43kA
DC/RkYkBLpTyLlh+LHwhrTycaeRoc/zM7Qk9Ot4qToFwB9o25ix5M7hXqMZceA4d
9zsqe3xTScwRpZBa3n+g9E7IIoUUALNcIxIKwwR+zABBZsUGs9Pl1nPKg+nrM7yj
CiEOLYQW7nPxi7TJ3CIm74ExdsThwOV3CzsXATPMpQCGvWEGSb5kSnl1mlkJ0KzG
2FS1p7dPYY5G7HxPVWGeYyLcif6k8Chtc6VaSVfe8guR0zxwaSbrtxf2yGr/+gRu
0VdMzCncCDUxfr7ZMqhr7oo/1Trf1vHyhrj4KooDZViyJ/xRhshkLq9qsHyUfqN7
eOWl20NY72Mc6KN2gOJinuV4ji9+g8/qyYi/hxCIN3ApVGQOU/F7lKar6gd1h+JX
WlCZHHDGac9m9MgOEqq9GtYSMPR4ZSOyYpL+eMJwj2pGE4ADKkgH6XpDYjSOvaKF
8Q+LXjfLMcl5nzC6tHqTYUtX32yrPi53vrHaJHl/Yw6PHGuJfaEHfPLPAMRSfzJJ
bwKzSorzQoMdCQ1KvMzp5sr2NZzi8bgpTIbaTusB7M2Pt4KbfUbhIpkpAt5wYxJi
WHK3D9oEoEl/y4bYGALF9QjyIVu3Zx3cq4eCDaYENLPlNA08bmeKqpOYp8m46tdK
Jh0aUgPCUy+uv/VDGPPMG6he0Z88glqyQ6JYHXwdXOERTJ6OvuJ9wucr6hNqvytV
xCzCdF5617eMAb05WhqliPXAzzrfKR/63rZ47aP5h7TAUaxk5O0rm1LFnydUb6cp
jEGb8Y1U2IoNhYDHRk04Gtv3l48OMzAg2y9skHVskgWLL81SZ/eaCU8ifc87uMY4
uxAKBC6BcsGs9qv780u6/INAK3S7ecg5qcUUz9fXebiaYPzdRRU3CyupJHW6MeQl
Zhgy9JPnD/4r8nEt8ff5ClU+t5dnCSWYxihoY1gO1Rqd1EU4lycDpu+FdRdrL10Q
ajyNxUqcYQmZnBVwr5+ozIxRaWuqp1ofDyEhdswiO6PtnpfTJDIdjdd+WuIOfAPZ
1m8hz40K23LHZ+tTUSP/Um5tkdC2xal3Ab9jlf9C4OZaprKDaZOhzsUoTsGABiaO
G4mBBDrb3cGh1sZ9SL3Jzl87Jf4sdjUjn43+RKQCZyVqDIHdk31J/in4koRipm6+
Ba3EGKvm03opxx2Zf072sKYTk02UcXCcWcj38QX4gVpJVBRB0U5dzpkxejOUkSUW
8squlJR3zOjP5XjgKV6oGIQ5NX5te41YiQKI0uT/rSP3vqIvkRbf1e9+yGSttZpf
FfijJpifZ1X7YeElZI2RJn1NTGrML5ZyqoXLEL0GFNMWS9+Yyd/YbeMB/6NPop+Y
R40EqzPkIZsRN6ErpOQ/XAzN9Ak+y8oai7PLPM88jHd5Jon5aaZCWt1qDtd7JY12
C2pG+FmLVceuRwLoyBvbgrJTNCTgpPXsTI18goNsZiQMjwn1uEYwDtB9zlHt3frI
q6vxNnxvI9eHth4pWLwcEWrFwZ73debVtRjZuxbx3vguT0dPnhO07E6ZyE/7SPQP
NretesK3BmcUvWgh0WIRKstO3WKcX/4dtdB83XHXyeuV1cEgZgd77vFHC7uW95wB
o06I8JMXNQDNh8K5sieWOvhvdoch1bLIXdGIgqWMBoGh1Rtrm64qzrHhh5YDMTZi
SgTu+t0k7ZBHKh2B8SWoqDX6p8k0MZ71M8nWwt8Vmv+89OvZvrqe4SDiGk6Y4Qv0
8hI0g515y4hMeL9/bJ+/nWUIi/bclbjWGkqKJlXz/sL7WQXWMQmfLTipX4bHMA78
3iXn99WSI5qmEuWIvg7kPYiGUE1GXFmV5bKkkLfQqefefvHRLwJo52/wDrwds+sq
rUnxAkb9lLED2mdNKUHW7aeN+iii29TOMJDe6Cwe5LFNh72PwWQ8zYWg9RNV/J18
zOmibhepQxoHcaeJZJ5K7B8dPMi1ja65pHwixoaXufzQSFufVow9Q6DfCQJ8gi6X
yleSRnSV6r8NwR9rXlbB1qsgbnw16uNAjOVEVdgh50+9eEn545aaNgFxy3W+C4Qr
+5A6cAGAyR6pgxn8NvAiJQfF900mTiYYGWcHtQCSfNTKF6YdN8demML3g25r2XhQ
RHdn7ohyaHB8k/5r5+4d9Pw9NNLqFP5seoqw+NIO7tvTbQk85V5NOlAe2zWEZH3Q
FBZHTOOshf0DOQ5aNaLKNAJ7vkUe9TAQ0lMvVMkdPO8O2KGpArjrZrNIpNqVGqF7
bIDPubCax76GSRZ4wCNHfTLm/OUmlBEUKHlooI3lu/vMgPPt2QA+xI4KXHg0FImO
QaA0PFaIDmQztiuQN3wimPHsQKXpm5vPVZf3kE4Sx04w3Y7+lHPUHDMJUyaLoDVl
Vty+hN5blvMo5MN/9VhNi48EPyQHPmMBC7/eAgJeFXr86fjmH2qtXMG2DKa/iArL
szD/Cfc5meRM2jPi5+ZQqh+cU/uFnR5EYXBiVOweaeqfs5vUArJnwWA0qZgrun5v
nYVb3zWCl9/FA3n8bDmVlsKSdMtdabXNUAlb/vffG0OwQmwF4lhuwhhFhx+z3Sb2
AQDKmyXhBGa35Q8+PPu0tTsrzpQRy/6wxvfCHdXkJk8xDaelMh1ITuP6HDJLpjcT
aN4Gl+Z2Q4pcJZdJv20nkxOPNdkHTnIhCkxLvCqEMDAutMt9sC3deteRiSobUHeL
Y6YNa7osyteEbUe749TxEkC9/lbAMRw6uzHDY1tSBnIBIAXp26S/h8BbD6sifMJC
2/2932/yNSlDRAnjxTdp9Rl2mdMOsk/MMH2MIB6umWHOVKXns3tJW/RL7jo+f6f2
xILhmYriDbnI/KXE6Dmrb/bU/OzCdCHkDbWe316NFvhrtXb0fd7UrbCuGV3/6Qkt
I4AkuMgB8ocWeiEWUUOpiTjOQLxYEGA5YA/goEzxS6/FkMAvNrcdjqf4O5I1ClB+
QqTLek95K5deTzlBlX/ci2YF9LdZ/ECkPvHYjI4KKdnEp/0KK2NvbrlI4eUR11TN
UfoGZJXrNYdrZssWB//JqaarYU8PUJ1FzLGMX8Tk0NVCXSMhrrRpftPN0pY7tJhV
SH+k7VQ5meo0GLG1M7e7GQ/OPdYitUNwwU1Wewv0x1CXurFXpKmtvshIYDvJ+Ngw
WNsnvyfDk+63ISa7Sz4nb9TUeR4oFdXREQWaxHlZJoNDdL+5Rv2DUlBcQJ0Zt/MS
31/L+V7JmaX+IX0TkEHnk59RysLtXUwLizUV8PRE0cOwsug4c8QqGWRK/65ttaWD
k5krAhlXHuItxVnJIt1WFEUVLuDqoBYTdwxMucxMMh1jPzq43PgA0UVVGITstf4W
5gINMRro/pN9UfWHTteqAt97TETnaB13ZDrLRrQ/AJ1Wov3IvRPzwojC0ahO+OPg
FAz/a4vHhlGwjLbrtzAkXY+Ro5WYGfiZxxK4Mu3+gA+iVqFH0GwtDG/5D7bmYdI0
qKIForrn+21Qu3KWFS7izDqGpvEiRCi6SHfzoTWB0ZgwyfTAaOIds9FgQ6AozvCB
oe63WkNXyglebNG2LZ+w4SPAikUCgncI4X8WxyxpGdLoLoVDlND2lqU7cqLpXu5F
9q5dAX8UOzeIPB4JruURtHCD/God0F7IypWBHx1J11wey6Zfl6H6esMVCxbEnvx3
zhbsZG2ZNDzsP4J8afg6se58A90eEGC/cncXqGIaoMbjfyW+FlqTeF0TP3s6zkzY
+vmOel5mKtoXjTPl9cvcxD0+Tu481geLNaxJnqXCraiGOX8UGUFhYyBL8VduB+6Q
tXoq8+gA8C2n8HwGd+zKBoyHs7bvFfe3ffnAE/dQa7T8lAY2dJZ6WfyiZOStpjYo
qo4iMdABS1QKnZ/1takGaKP8hoyokRVY81P10oJPC5x+ye99Ug20RFWJ1pB9uknI
wP+BM58czGEiZtIfCCWThFstylQZL1OLQ569m5FfmfSDq69NK4eCjKsazDMUAyec
TsShWtWub1XqdStyDk+gCnJvE9v3cZsv3hiDUEgRfacRjU8iMVYMtLzmkh7RYSdY
khNVIi46IF0Af8syXedGKUw4CcSgooSgHBPdZASENYr0EHQ0EunPlTdjcNhuJi7b
2STBUtzC3hQ6ceK5g0CiQ/UUiJ3S6QaszjzdrhgzcD9Rdys+MgfDTkrXGcWug1vd
8PQEVxp+cgWHk8gdd+gIgw/6lourXSgygGvafSvG07u7MCXD2i1l5pW2D/o7Z3j5
VGCqRGErQK64JJPAOl8Ty6Fd/gGQIYKIPQ1VWlJQsSiCo9PcoOkYCp3g32C7yv5O
qDyUnLYkXeMeVZuSEhfmMCSYv0HOhLnJBoqKdTo7Eo6W2jVr5rjqgaK/vubCf7O4
YElT/bojEcXZ8x+fWW93hJyaJKLuyNxlA4Dkji2LKsTc8htSzD1g6dhZvvKmYpwW
IZPfagHo4s/ug8X8r9xoenHN0d2l/7mxifcfVsXw71SVaKAN75IFIWMYZBI5Ea30
EmhyNu/NEKS4JnUu21Fj+D1Fy2yjCsPGjzN7OspjrQ5/s6PzpJz+WFfIooXs6hUP
aEmMDQMPCsSf/2SIwauG2nc42ERjyFJqx+Qj772qWEXgdRVMSzEoQ5e5hAFk/Tba
Y/WA/xPFqgWEspb6Y1L4BRcn9txyL1bEPDh7JENZ189Lg8l0/T75mUt4NjJ5lB8F
ZgDpDSEy/dsQCMXDl0SQGttm/PL5t0eApNGvm8YsgzDBgXc2pMuchUMGrqc9DTsM
ffgq8Q/2QP5BRu3fvrYNwWbKfdJrYhMsqxVSU4aGiMGHZKiRXEp6z5PmnpVUogwd
CdwELrdIq6tPGIgYQtV+hveiJ7/30D72Oz14LrS7SFOVVKwFOdIFq+Ag9Xbrs61n
kP+p+0wPYeBEBlcQRpxDGQheALUf5Dv8jRgFwCNWxg617Z588+LMwMGPuEDEbodY
UN7IUTcGFsnACfYWhVhjSyqMVnZeViIyWGhAGXsty1PiIk+AszRaGRqIZNxaJUr3
OxiKGD/ji4actfujf4XVvlZ0/YrtNA2SiWYURxg0WlcHTDcFumOVHwYaIj+17WXE
xrGFB8bByC6ugv+ZE96igh6PrNueqtFjISFFvwF8qbr7Z8XO+uKh3qGH+flZ25Xz
O6ZWHtrJxBpqmRfOpUqfAVnMjxkMIQeWHR1NovCu2g6lP57DPSSaxM2owmD7e9WA
q2gZvqOazyU0psGBmWefEElI/0waZZv/u9KVG2+jxYvl+ZBdzqsTofnkpq2BtEBk
brs5lqfvEmhKG/OeSg2gFq58XJerx2laLIFulHB5SjLyVqrUHhD3E8Sp0tTuGrro
TeGDpz7lRrFWxszStiWS29lq5rcH9/VH3iPHN9q2hLnpCYVJhrelT//jIf8JQmZR
DfQLjM4aY8ZkBW0IWgLngzjIZUk2jrzN7+bABss+cHAKK+a+XWMcnSiv1ho18RyI
KsHA/azn8KAL//ethKXAsCvlupMYuXcTH5SZycK8I/VRoc94KhFByt1zAQf/at16
xTOXErnFXJcBek5awVt6hM6ca5UsDZZuO4Nkvjqhi2ofBIul6JAI6L0sy+jWZXVH
mzU190GF7HZzw5veQs9VCAb/hmA2gP9X6OdsCUqasOc9M896EiFFRbzDOSPHs1zP
uNbdrOonG+jUfc6mqBdJ+q6vzZzeJuPbGnqcXBTMEN100PI5PJdAMFrhqvCUNO3M
7efTwuTC71FDSnvem594ZdFij6w+qf3gU2kmQCL/H6vb8IJ0vOuuXnw/CFwRiGKY
CX9Q+1PVYtDFeFUk7iZiHvI0R6WaXW7FmMWXWiOUmKxHK3CMDo4TzgHz/K74CBaV
+3tzWBKo1c4GR5x4L40gcMNE8aUL7xH6lWBTVE3u0sZAOutokk6hhk4K6BjKnyr3
8h4Q8CZAqYWRqsKJvTIV1pmE43mbegzcLbNp1Syk0QOsXqaL3WlU6oku/+NtljD6
YRTbEvTdYeSI2RjiRB9gXIr7dUhEw9wWgpQoHyzS51lGphFbnPlqbT865CsSWAsa
KWrHthUX6tncMM61tPulxrM7wLbLbRDdtzabKHiWJiv2brLk7TYeKV8ZfIP7MIys
MPXqDAcVYeKC+PKepPW1E85c7uQYxyvRydAhJLjXIAR7LkU6whP3QqJaaORMPHDj
fiXFKV7pOwgVgjeSl8aOTl4C1jhfNHF1vf2xRjmD6KOOHaAWYMhVitQJqCJaDT8X
Q6s7FnD0P/IKlGaBcWvgFGZzqFrPBdfc7GHenTspJRxDygINCvwkIPjqKZN2bPoD
GiYYtMtkHrW9yGysQ1wlvTXPIke69tgT63LKyX03y746ISufWVrLKafWWKwPVIsh
N7wFbyA2qGYHzHbh79fqL0MVnNH/68rjFf9EzsY95LQg8OlNTtM3iXN5UylbFxbY
AtuYCMWJvfRFJKmtciWKMJyRiTcneTnFoxLFOlGIc00j6CdCb+3hw4chBbzOjuw7
hlawUZX8C45rxtD2f38L8z7yD6OVt/ypoK5GpKxuZyTDs0JEJDYOjLiOIVbbTrft
9IXCd5sLZD8j3CjwVNmkGzewOhBOBdf4WQnCfHRy3R4Ydl4iK6SrfEzxSe0mVuQd
yMAUzGCdzMAusIK3bUtqx8RPWHTA5AcHtOJlXBanlPqwWM/t+LzmgDB1RtNrXW7z
vo0M56C4xBPgondDr1HhNio6CRYjXnlxX+TW3rKBONaHfrRfqNPhcS9dMTzXAEOA
0gUydQHYC4tVmIiIJfUIsmPmHZPAzk9fqQ4tQSDjtxm7afkQD+yei1ICOhu9dzj8
LkLq0QR/pmr9rW9S4Ogj1DWFlVOos166tN74er9bzYb5SFaQCxrQA5nWz61KTyjI
VvqPQPL9ViXIrGzXb9NXHdL0rIkgA+oGy69Uqj30ehrxUX5TnJnlvHT7awNpE050
1E0PBK09Txs/EEOJYufyac0evpj0VINfstx1+pQHhSb3/uB9Uw2+QJenObtGXtcu
fn8IGjlpbItv1BaOvAh2EK1IyVICBWmkseYr7/rB2ju6vibpTZuyejbXQnOp6ILR
xHj3oYW81fMZHafk+xMsSamHC73h0eVRjnD+cSmVxoXDC9W2Bljqb/h1IhUXKd+p
D480doVFfHnbFF3enhNTtBEEpzIT5r7cbWptPQ4EATtEAuPH44GFcqJHcA5AYohw
aXzcF9EI/sxqTanYTyOEr1UwuNdxf9pSHq9F6iaTiy1kOmLr4KCHN69cZkyKmiOE
HrstW1IYGkzQKGvHqq2CmdSNSAlUyO1LAkOWM6xr3EtTTsNOkjp8OF8eWq909uB9
ogjNB8ekqJGfybHAcOR2GM3P6HVL47QxAz8Hhpk0ZvTZwy3eASqULCqbckR7XUFo
ZWJG97jQ0i764UFfLnitvV90EYwf0gmmkun2Q0Jxw/DR1N6tBY+gbEaCGQLrceOx
AU0ynJLNcRA3s/1yKF358OaFLjBCeTpJRZoUZW//qhI/LqFRPSsTvJhrSMmFHIsC
PMFIUX4BTt/qG5YZO60udYeDYtbvjaeRBoHW6VKYwtFwe25qXGYkoFgN79wGAs65
W+/5J/znY+NCcYxjIRCdjceU9vgkR9/C4dJx7tM8Y74SNxvk1TYolaZxSEcWK2Hq
DTXaE9cXOnZ8xORTIxRbYYbmaXrfXK/H0UMbcEXIds/3aKV90P0I57CmC4zPR+wv
P5RD5Wyvvz54luCdODBNe5UxU65nvtNdUVPoXBhWK0igVaR3z63tObrdwHSkHnR6
FdADPb41MJrU+RsYPeb0zRsbpFs8dYEGqivFP5JvfCxfMARxY3lAvb3UOs07NSDq
c0EEAANfAwF19JAbJrbqSeDbgnRgadpu8fnDkIowxkkllmCf3dHMiFzHOEljfNVd
fifjnQ7GdtsseiQH6l3siCwHNUuYiTCN+mrJrodmcdIqMsPzzTG/fUPVjpvNIOyO
GXr+yAYTcZHBlw9wy+0rhKkLmE//h3/SvmYE3yoPZWoNMWjnePFldV3C49LBC7EV
oNF3atSk4ErJvf9bwfXht/HuzscgUv27Wsq0rY/cUX26WeHF4lZcP7AZfUDlDr0R
GC74SUfUidgNAO57sdAtRgR8IZKthjbHJ4Ga8r2aBkfPRVPsxEZw8hf46jfBlU+5
WfyxJkCh5nSYfBCquKvBFNUTNJg7cugqPawVPotwbnbz18t6D4umB30ToXoqq3Km
bVhLf+ImupLeDF/QvpaR5d8q8NrqhKpEjKwufM5StQbdjQSgHu30SI+3zK3Ptp+e
j5oYvQeKKPkBZcqv7BjQbG5swtB1hhCh4ie68pYqZMBhtWk8tpwEckxKKkuMLX/Y
PLRgX92KSz2PYnTNawvgu0Qxkc+IKXEVlKtkDNUy24Lc1U4TjN3MHMrgj34bcTIn
fHEhcjc+lKwHza3ii63TVR1Kq0ivocLmQ2mTTsqT9PHDr846ADjnIZY4zPwI02Nq
AeYRN43aepzcKhPTMQGxYLv7MhxLVdOgRaxaz44bBOGD9Jlu1AqjRRTiluAHYeeO
duyNtZ+jV8eVTwqHob4HAPAnMRT4YRiafLgvpklAsNugicBhSLN0DD7Wuq9Nj7nW
5fXBaqbTz17RkvnBNOhAAhL/OjRdLePleNuEc3o41ELAPSbaPPrDb4mFVsSa4+4l
4y+KrMihx/+UiX6NbFCjoPaWKnj4BpUQJ7KgLWLafMAj6ijLv1zLLeztG3GF3cnh
GakrVsjLR4SBjqoikFwIeaaKYOA/G3zBqrQwv6iMDWrdmpmrRSllPbKKo3+89ENL
2ECZ/7ZfeGYiQTX9TG22C1BalMoubzVgXdFVT86t7V72QS16o34pnw5pkT94slgD
mZsJNRzrKqZ4UX/t4QZ0sl/mXctZHQuXEVxY0ooqY+Hmv8G7pP+gf6LeOBKUDX91
dMdGooIIuexAyk9nsp1h8rovYexSpHuk8sIcJ8iQDo6uG1zR/waVjjP8TKa2eFvf
S5pmnBjDpd/cUd91aNmGNUu2rLcs3f/o+i0auS2Bn+weKbqv6iE2FfphhvKnAuML
LKm3yh02j2++s2bbl9OL3ASTqkAgf8aKw1Kagil9aoSFTD5i2w/djOCx7HNI0PjI
8g3iSnqqmzSw7+4qbWCtTpSw2/RFN5YXmPtInzSWEo0LnIFzoiPKbouorP6BPThJ
pCKA1r+94uESVIX9/L6xTjSmRvoW3MLu9zBD/YyvWdgflGMUowisHav/5hRvsHOQ
d1P47aDRMV59Kk1DvZ5bNhzMijdW1KdJjECcuxtdQFSqLfzfHZNkwrLJZTUk4aAv
0LK0kRwAiQyou6Jb1kwLWtQyTw6ZBWhoSAEtPpaeEcEKpV6AHzjRIqDfXFm/SuXy
AlyRzGTel3FD+ZGE/iG8vi0ZkxiF3BzRdb7RmcUhTw09SRg4tqmlDKqmznLmIs/L
Td/wY4MJBfIBzlgRc0nYJ0SkXKBl7x9Sd0y5r3n0PI3S6ZXBB4hkf9iAUWbEYta8
AnpbE6iQwuV9XKfzLqhLR7fSIq2trZtWvc5MpxrwV17Ymvp0Q6ZU9pvI73jQETbm
pc8xV2xlz9NCTohWkfSMRjGU0hSACmVfcloTuArHGulO56Wt/kbxTzYyFqXWVSv7
+pO7Aas6ZdjlVjyZBdpAzEXo5TJIX6ZKmFTPiY8RBMRVoolAdHDiKL7JK82HAmmU
N6ytC3PQejg909bf2jaAlL4Bib3pSJV+ZJOYNd7IpkbeHQTJFlNcHuEz3wpESqFP
+B/Kv415TMu/Tgs4eSJtrOgwhrukcMUw6KZRRUmkUTQ41krstOs/NjLfARgDqSr1
x9ShBvCoulvKW9R7JrsJeNIdHLmYNjNvVpqT5q0CpBKbiFPyl1apDXViFZ4ZsXGb
ZrVDg8cDr9c5FJXkroNMK/X9f9N1nNOotVMY/7Jb/c0XjzA8dX7Qu0SojHI6Ckro
n5sqQ9Bx+eB60WqH5uQ53LCpYNG30bbbt2LlcUtt4NcE7eK1c0EeXSaAT4fpiAaA
y6xqae0Ekcm4m1cb3rwyK3uC+afpcrhEUzUzhj0ZCLsYtqYHKtvZxVFCfVZnmblT
boQjGUXycgiMuTqF7hHRDFQ4PimN79YG+Zccj7JWlviXUj9eU2u+GNz1657fHIGO
ZA6mOgq0eKsBy6aDXovDUyKtjKZDqWcqV7n/9AyCWV+a0JkK48dezW84a8IOTyFj
7hgFRsSkr0CcUbJgy7tkSqeU7J1CI9Gfr3GjidLe1YSvDdYQ6Lq5Dw7+szxfaiYh
PgKo/WQttKT5+B243Lu5cT9VlYo6yYaN4FSmk3Lv5aKivLH6djpbjQ3eapUOizNl
naJVZ78w1+BwObTRv6TTMJaQBCN9LcNNad+RcSew8ANvuOCpcIxsNDGr1v5onezV
mSjRqewthbqvmt3c/svrUW3p3no4N+IubNAMIMbp1Bf0pBRF0ALA7nBTm2aGtWZD
L/lyUTrcdgGpLYHI8LcQ7byiYWhEVkDsJNzO819l76XboDtdBZrtfm6rwYvVzdzo
8719v7lzRuzaZOxAwd8055AIEDw1w9ddJWRB0bWxyMhj8SN5i5OlDNaPwp3GkJ69
Sx7FFZTK9odFXl+njOBeeFyjZ1iOduySwxkT2UUxxgDnlm4MF9yjw4eOxH03YiLa
yTmId/GMGPDkpcEBagqRi3+LhMu1AxbW14XjK0whPdyOwXRVJ2wBprdA+y693zwb
UfO339OjpYztd8TCFUGqCUMsS+6U5hL6JzEAJSXqBMA+33vzyJEtcNdUakMon9Sm
cYgggd3D4WY6JmrtDrVi1dqqHQ36NLvoH2832RdwAxw5ZvkuRlLKZ9sZjpFwdt++
4rpb6uWMCxikYX2Um1z3/L8QW4ME0ut3b0DSsjzD3IzglHY59qhtj5/wL5gyZTuw
u96GFBXc7mvNDTCm6t9y7ljz2rLZ8r9P0iibIejixCwV2jfUaypGVK7/ka2k64rK
6m8+kQUvO7bJGX/bCxwtr+roFnsw4mm+OG6Hmx9IQT1znug5ZVh0NzrDnZYmf4iN
FFBOBT8QK5xsQjaJwcX5jKn5trG80kdJp3ajkElJ4emeuyI2BQoZ5mtl6ek4awvv
fc/rS5QQUKGc+qOYYMAE4FNraTo3kH0e9PF323BAYplJc9WcDLZr88dqRDz6iJjp
TF1rmEmCdjUuV0R8JklW5Q3NIYDMMxyc4E8UHSAhYkY0vF7PLHrrSTPvLLYWd8r7
nx4LXMDpBrIZM6Zxodtj5BkQXCjQO7Av0s79yLaAvyojo5MXiQuyKZBtLBHzeH4+
Urz5jAHZkj1jRUpCW+/pul3kUAHsJ1YpoWinsmKBLBBr721uNcMXxAP3qALtQcVn
LXRPTRpP8cAtSU3YzTbP/uyRGc6BNMxX+UTHV5HSdoFqiP+sB41qiurWzZ5Ltx7E
yEjapgi8zbmPkycsaa5tqu7goJLSPoT6lotlKV7CGLI9LBXHQN9sXbR9s1SSiSPD
Me1JU6X8U2MLu3RnoAeUWwbECtrffRr2DwhivfdkUBm3OIhUuMNKfKl08QIoeZ8l
R0tqmfA2m89VfRNnsSeGI3xmJHfp1xU+3DqNOHvClZoAgxp7W4B2skMosLRvJwE+
U8UUBqjSLYVvAFICvrNBoER6uHzoaq/74SJR8HBYL/dhHFp2rsO6BqMFC5MY0qlO
cPAYx5aFz/uKTHq1hvAt2BZaJsJsMg8C8uqozfH2Y18Yiv25m+fRVLJesE8pkYs+
3MsM8e1OGExkGMLrCtsaDnVbaea/smV/sLD+HXKDSCavVyg6i+aJHZMKTD08xscj
5zp3YgqCsEMFog8fMV9i5fh3L1XhpNOvcZfJ1XQD9mH6XhDI+Oibmr6gYkdh/aO+
84UoUqHIB+uHXbWAp2cpejt6/pIjdlS3xIDbs4cDw4qJY5hnSV7xH1aKFe5nci/j
mLylPn+bmhw3EOfYeNBHcjKh0J1erx87+BGXkd9lNq2bQ1v2FO813NxoYa+WXowZ
gV+Srdn4mHbwhq4SlRi5B8SaxC4Bkr/yrr40Kxgb/zfXu+WSY1wFqU7NhwHd3mss
tP1TCzA0yalCVzzXVk66lfDOZWQAnzPLgSq8EZdzvL2168ibmOLWrecsu54oUxdB
2baW1/hDSKk5jSdk2tlq9nIs3fNkAREosXFxOryYLnj+RYbVjdymIRPmENkO5Qph
CeL3pqAf1fq6Jxj0RMK4eulKC2YyczACp8Q1D24R1Su/4G/E5OlezEC6kBRyh/ry
FTLGw/ipjb+fW5UUSw3z+Xv1Cb6h3KxaVjRi1WeLHiVZhnxyuYD0896tagXp15zu
52vjc67gXsipHJjHDsbz5QJgRHn/3I9qzBIbtRWVYVPLDxIWXo+5PeU7m1mQ3eUw
1DxR3OP0exlF/3UvA5SF4uFsHjGhpuywPTEYEKDD5aP3d4Ak+4H8A7TdXc95hnm+
jUVTV/da4mbY+rZcU3rbku2MG4VbmODVaalBnUf3WCxQSJmFYYIhgK5CjRMu+2hI
tFMa43mO7+soMIUDqpJQPjWD6ZeIug6hUBIxHuPVaqRAKlStVFMNwI+EjeSoV0Vn
VaiPqUxXtlLtqv2QdetYzSiKT8Art63oNjs1KmyzOO8HSI26XubW5dK+7OSMLdOT
jrSRJUKo3hwmRPoDbsA5LiWMMb2oKq8tml7LhYJVQeSSAGVTHWQ1H5XENZ66q2SX
rTfv9lWXFcAxnbz+ptw3sFhspVg+FnVCKHZdqKFpmkcnmFLBUFc+/G/jJT5jqiVB
MMh0vUJ6y0goaC6+onHo8vrso6AtOiO9My/Yh2IVoO896v+XChd5FATSwqNuPA/Y
4jjBva8oIoEdFFL0Ls2SV8eZ9cjPiklbWspa4wg7KFE9s3OOp+mjxTrojfips6G4
YtzBdqVWaVn9JduZKryvEIjMM0v2wQ1k1ufObsAYEPWLKvew48bube6FZ5EBmfTE
0T/PdIKpBg3QmLMyMAFJP8DExlMWzf9wxtpd5X6hGf5tBhmLkjO197tptxJNtORU
ZMn1chJb3ZgS/yi3JB9EUUp+NEHpBHUI+H46+R+zRueSkGeEcDhldpZWo3FJABBr
czTJwH6NeFYD4EjenWAtowP18fkkTm97mkitaytAS//iEzxjITokR0BDFXJ9HuXF
LQFcO63QVGjlBegCtEQpUcBClsm814MEH2kOPg/7l+eoSqQPq4jali6QVRtbMrz/
ZXPpi9bWfReWyVtymnYXfdwdLjM+DcZoTO9lXfbSN6qoLi91ucaagpDCAZmacnpV
d6nMhjMJ64rsE9fEazqftm/K90kPQY0tWV4etyxDyTbwUEGESkelngn0qcd1ACLJ
m9knJ4fNoDRCgDusuiwqOVh7+SKq17FI6jWW17i0ob5PpLiXR7u5ImiQUL2z/Nnq
Yoo7WPULwm7Owef+ceC8NdfgcY37XP/BpG36jUlLcoy9MQw1ZKdX1ATm4BO5VF0E
WH1/7GECIamWu6t4WcxEXXLZVobwQvVjC7Mg/AgvkAq2HkYffWsUf6IAGgN1yRPv
OK/u9gQobIbx3y3R/agys3bXReuxjTIqd9qsGicuSNSTq5R6rW01H4R7ebylhl7o
PuIMNZ61nuDReOKw3ka1ZFXjadOMPX0iIeRm9BRmLuGhfhnYMxZmgkbh6B/9PrPN
2tcsisHwYBTi1VXFVHz8PwQBUbGOpUOlQ+nEbpS06ryR0ZS0rGKLm+nYsEF/eKpU
o+VGlZeNWaXtURh2oG9N27f861PwNsOSq9HZSAot1I9ruguGe8QeFlPKJSJzQIJP
jxnJSWmRrWRw5piwDMUtbEepi8SsIV2g5Nq9jlxOtl+8zujvBe/+elat+7lkvQcO
ciFUFh7NjH/G4AlUzlutymp5tnRMWM5SIkopGr8O3ctGRrd1U5V3AanWv7v7gSVy
hVKGBP4Z9YPEG3PMN3S1q7sKbSjzQi5R86SNEJFU8KYpDM5VKPmhi8kUqaBcthZP
SffYb8E/Ca9I5jXedjH+AmgrmEYL6c9httaQaQNCrle6N2UQKxJ3DYAyUH9a/rUr
R9JkNbXX2QW1daZ2W229h3HWf+U9D3OHLeSdUhCWfhn8bd2G4KsKZzQGs07H/D+G
AizratdvmYzr1Hv7WvkbdGQR6NBcitTDKP/AMFgX2hpngWSWNX1I1G07dYA1FCVM
hT6IxfVgTu0LNapBlqi4vYB7o9oM5jaiZjy2GqTt/48pxu3fXpUzZbx2HACBUUQ+
N98z/EJWzzGjekXK8nJLpIQLnkFrmyaXC2UZK1Wb5DhHn7E20TD+9BEoZwQOVh4P
SktgN7fr+X7O7LXWHX6JPwjHeAPvzCDlZtHQunMGm/ttkK4MYRdOcT62t4mI1HFw
Zwxdj8WfzTvozcB9UiAIUocilHtxwYsmqjC15+tzI1TGctrtOs/tzNKhud3xqzJC
l0m5rRG8iPRtyKI7upBiUdGVsgC5HinGc8Imsa8lRHFzMB3RLY3zyq0JRzPhY9zQ
PVoN4IpRa/jJxrrQzdykuoIgY7R249Ga0qURWxSFvzgQ28CINP5QyT4BhsB9aeUS
prAnwDqccBJAQuSsEF/pzTY3pU2wGKLaMQH5cTeHFtVYujsi3+UgB44gYMHNxEzt
irdCjH7lf/2q+U3ytr7F01BxY+ArH3D25EC37ShOnp209VbO9LzmIp1VDTuEBeop
2GXWdPsjqYZ7+lbDfzNLp6Jhe3q86vIfG4zseuzcXADtL9nmlgCYIKq4hOqoomrG
xKBvvmQHoCYWswJjkiXeFIeZd8ojP+xX537nCbGuTXULgHOZYZqSJtxwbk97I2cn
re+HEFmRdhq+dTEqnLYklgtxfkZQb9VywzpJymyPpqszYqZqBNaVFj3c+ljTbpWb
/p8gWCkT/XRVRrtgpFGPBOx5Ekk1lh7B9juViBuh6OAo9hCzSINxu8cuWlcEfrtG
GbCHbd5HNqH8y9yn0gObxjo+uvlVYSiewcIgkKfpvmBU6zD/AsEwUuwWLHWmzW5N
gf1kjC9OSZKAtNary1DKJm33RW+VSGOHyFnJ2GGkJWOMPoxKtA6o/l28c7jT76iv
dY95fp2Y6fvFSEIUUr3kL6hm3aRwdlsFSOwbcam93dD0NynS5cZvJCl82io38yB0
rsp+p485vCE9t5Rq0KzGbLA/YYG7DsD+s/rxdo7N1mPnjGY5W9EcOS06AizCuiAP
b4ZUQwwBVhJwHHHnJVIfAkpDRhmBche+85YFQv0eJJ2eDSYNJnQNBap/nvu45Vq9
33FnJMeUYKeodIKN7UKhuY5aCyDgHoZmcRmI8JwCKXIEw4+AAjhNqOCamLcisJeR
H35xyeRpLgBRSfCfGN22W72jZT2dWcAs6DaxOae+M5m4PqwdFRzh2PNA0AZCELpZ
SgjaB8gmPLQZGZMdmH7V/45OWNzLiCitD/Ia6F8cdmnmfOZfhjRjHAiNSd/cj7+d
8H9pzoqiJwahTGvjgfK943NbHMjTp5ue5FOxbCPbnkdWavzdpGTD9KqK6xXt5JRi
7rJIIWdM53fBa+gsoeDsnaX7C96lgh2ASDZSciLXC98f7Qq1xdGOMCBFsCo6Kyiq
wftxxtxQlfbZFExi41eAbZlmmR1ZPhD+vs0BFdqSmI3hJbD9ff9+Lk1J+01UUjgs
YX98xjVLk9m8Ao28ntvnhVAlUXajG1uq9EF/3E09MxnFSbY47oGVj9j1MaPMVhpt
FE1HiSDVNE443/4fso7eQL/Zbdw+eXEN3nmiXK5NAnFNFLOUzcDIWQw1OHiZjKLB
sGMCxOlkEFHdVK4s+mUvEdd46y87FpNwFlXN5nyh8GzcvcxzY/QE66N8phq3KSZs
6M3ZaxF10OKCZLzXm8/YSN8Tv7DcfEp3UnaeCT+Okg/JARhs5bO584AxJI9KjQOf
aEvrmVaTwB1GNbkNR4vWrVObqMI8GHv6Z0b8kMjcmkCW5ylFXAPyTLrE0mAAa12Q
vmAF+5pdD26CWwQrfPo75s2Kg6LMpL5iP7vmh9yfo6IUAfJc4JSTklxwupYTh8lk
xdGQKKH3OTtW22d3eIlE5nhnMnv3dO8uiZ2LSTgVMD40XbDOJ/9D4dDjQqm8pzdQ
XwV51dzY6X1L81lscjQgEdq5kWCCl8gDvg/VFVvCXWpVotPFAjAUA938vI3K7YQV
cPMp8AaG+aa2dH+QFmTQcdZOl86P/61ZjbfOuiE7vfRJWBiTmBbh0izGV+Zk+lT9
0S5CO+wtSfCDYrwmHG18/1Dt4DLSgRGs8Q7p2PPsedqYlCjVHtKGCeHVbIQgylQr
HixIOrz6qRgkvraf9w5dJgUBvGGikZiWc+dsfx80jlpPS+jKMD/+XulXHpz/vfOD
IKowYteW9JiBUFNZaGLI9LSx0pP/zkfdYm44MlpZuV2xMs4ycuqd8irFI375ili0
tWjtRPM2EAoXhGfJxtDR12zcdVW8h97x5ToUmco63ew/J5Uvn7l3v4a4sHOCf4t7
FntrmscjFyrDeNMpG6vzeh88aLCm9uJCHtcGAM6NzuxJjT1GMY7hzzfmLGkT7tra
ximINGYqjWNIBHN1zYQNQZAsJ/SB+9vWAqGrO2fbJqMPaQe+S6w3uzGwaRNcjLGV
FE76erXHWdaU9pV33LIHYjtCj9GnaAy5czr5KtkACPaXrlFedqZ7pk6RFecpCdX0
2SH4tlGPMo7hwQtnqxMOLegIAshLJ/QDp+iqoQRsSKFKY7fLdK0O8Cv0JkZ1ZKXb
Xi4kNSWS6LqpRHtu6rP0IAzP6+Yk6cuKoXGiDrNurR3jts13zfUzitlFpBEf0bze
vXgUNi4+W2uPzI0Lfhu5pBT4khTMU79sjhvOAqyokJDk2f/Yaf0sA6UgQ7c4hHTW
vLOTl5tuOBaq66jP2K6FnJooY95+YI1kwui8So3SAoSPJ85rPI6CLYbzVJxKzes9
ljaDiYEou7/Em5IDZR5CGMFkEGUTdK+QLzytAYq7DtHReZrhPa+RQua8+7kJ4vCx
osN4QMWDXqZETUZRKAA43GlOC/DSZgY5qIX3OUL9VRNolOIPkCsVq8/697wDIIZW
/NveyNr20e45IqMdee+4jq9Ghsl/ZLE4iV9roOkqvsLQcAvWSjd3OlC+oz1vs/C5
EzkFR1mbGwM9vhZH/r24mCSw1L6fxHkS+rstv+iCXWngPxe3J8F0Kej47Y3TIpeN
QzaucSUds2DxOXHcwmZMrZ8NPtTYmzXnN/SsVGeigOUHJUkxQNdcCh1DdnLzNv31
9PzxGkFPfOfwqe8SWhfoN0q1pI9e4/VGaSJebQCwZDVZGGgBcrk1L8LpRzQCQNJj
7TpDQIcr0F6tOwlWzlMsemSUVRTHoAYVLl7/+57Anim/RhvicJyoxDjnNYTPT1Bu
cBP5bfX7/38Kl8RoiCf7f1RokrCu4fqiPaIPY/WVxEy6UgcC7a44rv+xY5dkg5Fd
Tw8KVtIt6lUFuUfJNxm6shvlREuT4YWTUP1bIBfFIAeqip2ShBzEUczu7ARoOE6t
VFFVqbyNfFnCD+RhopJi7TnZ78b52F6vSoVKP44xpNrvx5PCR5kjb6LQV7sTTMfo
E6GYrGQE3JHWDVHH8P/N5X+feFYiD1TFDP3IDAXxm2XQIUCXbiumFc+QnFXedeSh
+JUL95bZlhfYLPb+d9DJryPL1wNe3XS0N2Zpk4VMqXyoezOYd1TBD/sjE7u3TmZy
04nqL2Hpz3p2r1O1XJM5RI+HoBBgKrGmeyYXv1bVqTn+VrjYaPcqUymtH1N5gYU5
owwQ8pC7a9vRZhf28jKid6No8eYRZ55Zuz1Ax8EPgCuOO8GbslPYUHw4U2gpgLvc
4RFzEUfE8AKdbatYMY1F9QaP1mQScR+MlnEJWgVptAscQvUgHZisARJfVsvkSLab
3XcNzeSCxe1hZ1YvdnANDA1dSiazJmtwUyBoYOi+MZsnEf0vZwY5GXV3qvrXnfCg
0TnvTHB1DkgiYRZ0z+j4ji0pptJFw4rofJQi8eiOJVEm8zz6D9uMEGbd1KgUFHfm
pDMbBhtJqtrBGqffR1un6CC29PWrWptQWxUQsnc7J28jxzje2KtvCDUt7tg8nmYc
eAsLX+peIX62w0ap6U8P5mb7ugE1PTqqbKgtUSUJ71FI0vhKXFmvb4iku70w4NcQ
IwvzQbOVzQ50gNLax7pujGCgkBVpzSLoVTmeuGQ6zV/fQMDn7iCLGvsuRXrCSYX2
pZP3HpegXXvmb94nF6OyTAsv1sA3zURGDMBTJQ4DxDVU+1Z0AEga/ryzbqyaeSmB
OYkCekNtbw2n5aGw9vy5Xllke5KELKqRrhE6EMhuU4FNC1apUOfPj4eQMe6+Lb3j
cupvgj9DdcGQIOQ3eUPhulGkzJsoUmd+/quLn0SnKbNEetWFK2ubSMsIWDwUuSwa
yTW673c4Wp/nMtqKMV23SJGUzPU1R1cIejz0mdqkDj2jQMYQ+jH+3PRPwyihHuCn
isb+vfAxUU0fCbBktaeDRIWQsDGbJUtZp2K8BYUoyFmov5543SK9Rpg+X9Bmr5Jt
ccNOJRC2bRf+LN9Ohv1wfYGcg1fSmDZHBp8xeOsH48+LpwdeSdLLNJ1JV5M+E9nN
kdk7cMc9/0c1kTX0UFStaUJn1l04zSLn48QDHL4HGgaOKIHC63wQ+NInLa8hk8c3
n1cZPqDzLMWdmug+upHD1c2IUBoszhVoaYO/RwNyb2OhKh6qALbmrc6U6OHKLDJN
ZxpDbX6oU9lc+2241MMUsd/abGg8+rYhcBWBiqeberqPyPNee1HzOQSgyIAG0wEL
rp0qkpFe0ol+nsPIcTdaMLaq1kv2KMJXfIX8RZxCBRYMKx9JcZmugU9Faiw7aoB2
PLcghbV6OoUoWqDmZJZM/QIU+bZCVrtzipduU5pCAiFl+kWlws3u3V4B/7J2th3j
NzyE5F3PnGQ3XprLXZwbt8vw749PA6DhuazqZfIvBx/vTRybZyuwyRQESTeWT4rF
aRf2CvnVxRUMS+oDwfw8rMuJVZsjMPWX91m7jaiBcqrYfLSRgBTMWdl2tkUB94Bt
tox9cX0f2S07nY5Orv+UC1P/Wp7/yMeovGkhFgx5gYfOacba2d+7PZ4l7vkug0YP
OBFPB/8dzoEmcbdxEXVUEUw8L640sFHKFtdb+dnQ+j8p3ov92sNAIqtX2UjhZ+2z
HrCozGlrkQ5Mllgqnl8vxdmCc2QD2AvOsfDdID875WJAbRR6fF2VTb0gHuo0WekB
4W2mHI4szJVtNqaV8XUb/S7H9C01CpbYWPpavuAi17qrV8NTGbKZhm8eMuqkgOEW
i+K29SFuYIUqDrASCcURSTkHYWiaSh81lFhIgqSDE5pT1C0kxOx/GiD93CfSA5w0
H8QB8SNHoSgo9H2JUOxf8AC2EFaWLKAoub7Z2bdau+ISwJZmEdbw+YX3KB5XNGfp
BIqiwE0z1QAEl+ADmEiZQ0sJ4tRwp6+AHGYXWuVjONmYCOdTQQC1gXgKh9HUnqzU
cV9bGFX3/46Ax8aqMRuNpLOhB/P7anv/kTQt5cG5zBCSNDiZS8ObVEIP0w7K5QlM
DG4phEOoGhoUpTL+nUiGkAG30v55KcmDGH1l9pj6sEc1zhUBBdT9LjZdcxKpRf3K
1qihH/8+hwEtkmA34LcF9RvmlZQi+BEu04Ely6MY7YaG+kG7aWeYkUc08HzgJU3J
oHPXyKZMYgs6ghr3BGdIzlll85TYxmz6YUv6eyEjFA194YvvbNUgj1dnoLfX98j3
PbDcKWI+mv90CS4iosvs1v0VE7cOU+fEtd6XFqgdmz2PDo3nFpFHiQJZ09BIDZkn
YoPjYPrzDCs2ljxnYDjGOvQDjso9fCFx2vYmX8dRUiesGukcnhTKKJQG6nNzmzV1
KNNQMnqzkhK1A4uETXJfBh0/VRHCgnC6CJsNKHCIhf/81WZAdSL9LPu6ZbsHTvbk
XGrg70i1nuTGeW/DBVR18R3jMTQ/vCf3w0SbXfQKfcKg5TpJIyPTc+wtwGbpaWWY
KvEAJ60H/lGvynGqCcBNBWJyffQYmIpYMILqR1zEyepOFgD0esa55G8innJyU/SK
cH6+aQOM05/DyjznsXMlnCbaqVHkDfTG7VFC8DGp4Kt+y2qm/qzeunOkDd7iRQHr
gnxHjzTGYyJCVQ49wAMEPU+6qV5QWFJvUunkv7/AE6HQHP5JfdaFf5f94T+vHnYb
Oya8iks0ieNooJS7vbeudEk9BtIOmKwmtxLSLVfGnN3SM8ZpRZZQx5Y6FdKtDGRm
Db8RF7vdFrZ9SWnH5IB+00NkY/czCHZi3kpfCPijexVFM+mxfaw58+k5XdmAcp4M
+pIEvoXM5W9p/dU/44cQ68hvZ9PTpaDtKTsH3YUUb/u4fl3s8Z45NGw2XTjOoFg8
uzLTojGKT+NwvsB3I3PVJYVUwAGZb80ZeBEV8mdaDbe11FjFuT2X3hIQxOnQ9MaQ
zIxM3eKRKDZc5zRD6jIUAaX+yhvAat0xVgZgDN7QpvEOr7m0ysYI+spHgPr4LCL8
lbuGjoqQ/yU1c/eEBLdR+EzB146G+qoUrH1sc7Q6FrdWDJR4rTulB4+5yEjWHfDa
hdVj8EF1/z+9VNeqx9v2kcwUH6U2EHNRqEybWHdXvx88b/k8CATLkUQU2cgGm+Dl
CeQULyhQrMIdFv4l2uHf+tBUo+DTeoU1Azlt0sg9G9CJgHQWD77xYCjoO8f555eJ
Zz4euYHK+ms5l5H5nyxlT3/SEeGVXfoANYJQqw0ZbR+Pg/4w/msucZSXwkKaCT6z
eQi5n+wm4+Y5Sv+YodEi/kndLSkS9R1QtA9guN7kdBz0yO806FMPdITxmZF0n4li
7wY7b9dXKXPNG4+6Ggh/U4HiIAb0oQ4YTrTc84PS1ZVhLW2AgFyq2yCGPRbL/J9G
NT/IweiUIs+ZX2KusLvYlgSdtSIvVp47r6day2wMeyhPHxSVIT709kQv4YeHMrBs
Mf8m7z26mdCYXlbMI/btWxVnCDaKxKXIHS9A5LjpRuT/rXcUBJLvrdYPGFALwes6
9FUlUytnKuoogzsytmyEKmzD7tmanENODAq6Qo2sGvv3axX4dRtne6mubSJ+ywqR
FT8gn9tBmHUwAHMclUaBR70ufDoR7234QZ9x243peF1eOxqh5wRvyIw+wrXmeVgM
kp+3wwsExh3KJv0iD9HuENpuULnMhzgRY2jxp+lEz8aFJN2y0+br8GXdlftZXPNx
D0IZ/f0hlOb09I6KKVijTUzwVUxyL2RfYHVTEStvVKvZXLvLOgb70WXSw7qMZorx
ErVGoP2OBZYscZLtuqCkaGWI+OmrJ+j0eyMj1EhVGnbWRz3nUmmO3wadRF8YmN3J
6K+pBAAu0vHGePhXZ1E1yg+DOYv+4IRVU9ONMJh0WjtRp3uDYTjcuOM0NKroiG2T
lBGDdzbbSuJ2h9kUAkTg1EtXYwkvLheDYl9NsYiU/wabfCiKEjfIZ7UcZu8zYt8m
c082ufBT8TnyJhRXMbSegfVQKQRU+nu3Wveki8iXFzSdN+g3yZgOsjAgio0Uw36t
sWgUxOFziP0Bwn8mQSyci6b3EF1Jr7fYjDr6NO87s48sisnB1aqf6Ne3BbXIx/Qi
84mUUNgQv5fw9K8sAAl0YTAw1EZGOBRv6sbNc38c+E92JpcUcf4uL8KOpDQUjeVU
k2HNNRz24wGBL6s5EhGc4j9gOahaIldIXqhi+rXI/MevTl7JDgRdLPCZ8xPGdcne
OGC/dFZco4fA1LIRW75XYIof5z/VmCMx+pUw73DEItrvEKciyYQwTbdyjnME7h/3
IJoSu2zxPFN+VaAmpF0X2PQxFKwqS55wCZRIVJuyiKQkdddLUGWevozboUFvM/gG
+bb0MKGEeWKnxaVoRyRkOsLIdEGurxlwZEluJ5habyfTOFnVVQlh1IPhpcCRsUwV
S50gvDe+Yk6cJMSZjTcE7g0xG5vftdd1DodDPw5t3UwB3NOoks4kyMWOzHasZH2S
BMdA+d1jSzzbh1fQ9HMEGGyTUI0v5FXmpCOT/QR2O6qt+XavjSVz1IYVHZjnlTLh
TaL98XnPZlFa+qcjkbNmZfBD0YyfKtGuB6RhcMTvp24IOiCMFd3jGWWKhS4V5kip
PMA7MyJWcqnMaLRAzgyLp0rZ8CBoQ++hDqtwI724Y5qlV0DL3taK3tx1he40+euM
hKSryk9/rrnBvC+jTr/I2YSjsxznTCV84ECK/5ZYncewdbADvyIoQ1ymcaCTxEUL
D6i2RPBPrt9AE2tXcrLUOVxyzO3/En+pazJXyJBsKSjjC/xIDhvEqnm6WahDweSa
DVPCQ0Dn0vvv4eCyUWLJbc2ZPjyt0IYS21ZgH5z9E2AwlF5BjxvsBUaiS99mUGGd
x8lRmb6S58ViZKCfGyA+A43Om4nmHZxJLD0ahxoBnk5Y+4vYZ7Wf7NZeVsBOdWc6
HP2YfV/jqzChYdAVgQI9xhvcrkPNWFizolrhu6drXMTEwLUrcsbY9uVb/kXH1KtO
Eier3eyt6a9vbm9V7gcLLuDmIK2ceVOKXkdOqpwgX8/fCXX96eNK3gosiwI34JJf
dLe4YYPStSu8HGhp3DGCa9uAf+vuRPvGIvmPPXj2HWAfgQxEwa5fmjZ49yWIl/F5
pqGclo8mNfXZW5UMMHyHRqb+J4xbVkr/s+yBj7+x91n3/olG+S6WBzEKpZHcnw4F
xi0+EwKXODRC0xYuEWrXUgtY+Vn4JsP5vEMi/uZay+zx0NpFwSMVv4XWgU7lIuWU
oQWOajVZQ89DsWnJUyRz+bv0a6Kg94Xym1soQK+p08jUhmuGx/gdeVWAADKBUiO8
uB/6Za8JwGRYimopcW0vij1mvJlq2yd8/mNJ7sUISNRMXj+JJD5jSDyH/KDrljaa
Yh6zagIixyC9maGyNUeBvF6e0kcBAcrQiHk9yNLk0popgD77zC23RLZz5/hhaITq
8TcZYv+TEgTNpsmCX23H/+7uPE9S5/Ns5bX+3SIckDnNCoq8MfShwiP0bSi4MNA8
wFBrCARS6TwV0TfQRxgohy6C2rlAgmKTA0XlBFbh7oZEf0sQNl2solLFT+KjxoOC
WXCY2ZZNUv+jwbJHlmrWTyqv9jdRMrUPC+iuUlkwCdRlHk+i+SlGIjoCPXjuoROB
Yo0lDBr3/rkyjTw6Gsrz7WnCslflv3tJRUwdpuwoBMUe7mpg5x/WFPBVJchcK5UT
byarBSqSU+71xgV8lgWloyCAb6GrImWdF4gG97CQzE/1nsWmrdfshp2Nm7N5lGis
h/jMbMuKfi12SUDk81DM/nv9dTPtfbFLMz0AwpQ0yLZ5UwepuWjaJD0LrxDQNQe1
4K4O1dlI0x5pTY3VSZgAR4MblDwX5NmM+rTySMlxztm9b7fPdnE8btphnOEnCPvl
6ICoaZmNgiuaPmPIbU/RUafaxP2Ks+Aeo4RapxpEUeANPJv8cTJGRyIQtqlqm0IC
6h/OqDDDfNkRafkaBDMBh0M5s2a1jf7t1yRJnZRGO3+4uyNbJtwu2edfHOuIfyoj
BRGwuAV390vyhv1BgYslK8OPnlPurOBQwKG9UZH2Imbw0r1oWwlXeqavQFAp06Po
uJ49/FoUbTtXFMmLfprhUDKMO2VGA2K1/GAsSyN+VDyzW5j69rxyX29fIO5cFrIC
VmeadGUdMjLYNDM3l51NHytk4JiK1J8D91g1A7FLXvC1ty3KKrHac/+HK3jV4Lvq
Srlx1Hxak3i1uWAGNh8xN7GhADqCB5lRqDi6u/Zukdjkjb+X2EFULecg340Nk8Me
7I1UHGmtifBjYSX97y1EXz5IS2Xiz9PnpLsSFf08JjAk7dHMgRo4bGdIDS/BbxvY
gGsMTmeZ81Ia8aeUJ4g7KAzvSpyppwypsjIGmgxTe63mD3qbdRIZhXxsYaFHuVBR
WC8onTcZWvRUGvjMmlUv8WkmUyCBb51g6hAdvijvvSVS2nuzloIakFmnJnp25Iza
Vn6p8W/pYcKlflmkKe47aIw2DDTclXhAEDO7XTr5CpfZbSkl3e3AoZhi9Qx/6upY
McStPuYmZ5HuT2lP5RfyRKAp3o7u5G+JEqjb8HYqsCrPagp+5xEzeEWsw/KJQGAs
fe2gB6VSxrI2lkzqKRsgioyeTaaXA9QgKIPXW5erFSexg3+FHkxOBigzs0J8/LkV
Quigplc0+R2FnUv1lkoyivA51hQhKDL+n5uTrLSyZNUdb2thf5dtnR9jerdn9qad
rheOwH8ZKCHHXNn2QR4dkyDEm9d29zbXmkIhkoo31Q6ljBPilQtZlwIvCvGt0LaR
ge8VK8WcWVgdUxhQjJMRuQovnoaKYql7QnfsRBCxJc3l0XpZsp2TSzQ5oWcJ/IIg
g9drRQ1Yw3o4kXvu+RSKNuRvFWi2m5GkCDaR6TF31uB5+BZ1UTQpA6oEvGax8u8J
GHf1de540+5a0Jvh+JbECiHETRE/xBME2Tvmy0qEKwZI4fmszUUTwGYh5Vkc2Akb
XhYqanpRugQk+ar3cx8P5DCZjyRA/4jJSeI7VotwFHuCxxFRFPXkIYOheuLW4pv2
QbiLqdN+biNV9miKEiGGAplx9O7CEemOBPPgLzzYv7XK7woEdhCluKbw5q30BoTG
ZmrvYjubEAm1JKjZOqkvDTUfGP9IAzubxeN9LXneQ20rGPwVnHD5rT+2ghI9+z9K
A6SsWGuBssonI0zagJxzYtlwRfgSBQlu/BT0WBOR5rZdIwUapAtcaGX7r61uCZw5
bLRsBbUflrRIKOxVTwtWgAJubxAKUrYMxRC93FMmdbccg39W498JT1YkuNq5AmQu
3B8cHfgCc6nGU87sIoZN4MIoNhRjOtzSMxtotuVIouP+QiNm81Lhjk4sjSiZisFq
94YZEsDk8cCEkVENbS/1L9ZMVoOpfMJZyFMrYBnaKnPmlZLEVUtsTJrFy0Yy4qz1
cePr8ch41Zru5iDBmg4dNyxPxUk4bFxjdaDjLC4Wvt4Sf9HKSagpVfcicpehnarO
6GiRzDzU/KzYqTO4GMvnQlSnZp8KUDj04lgPHdD69hbfz2MSf8KHuQtZyrhzGExK
EuAFAduFqe0vW5tBGb19QzfwO/UsdyQkOxvo2b6PjKvFWoxKJQHWkCwYpTy2R69K
HcJBDnOSsv0/4NjrIwhPvdXIvUI8S01fmv3i4BSQjCHWKzYQ4T5sCWLblT85YW9N
aaBriACpA1sg8oXJEQcwvaIK6avtFfNB0FR7XyHGq1FFUIfq6tNbZYz1HVqhePVP
o6YcgDf+qDqhUc5fHQknKReFD0ahGMdkijxIJAkP/NxuKL+F1rDC1iu3qMs7B1RW
awQkFZe9fdPJUXm4ksRibmy+ut1V9IbL+qaPrY4tWexZDYD4RuLj/tVehFWL7ibr
IvTj5IRcM13ZXbPpkSTLGPjw6L0OtQe9IDGjDQTSDH06XNissLEFd2w4QTqGetHA
SbSzlyRYpvybzUlzpNJUpf96Vvejs4MHhY9XmpYp+juwplzEUG1SbG718oEHUu5G
5xPTp1DjXg8rsLsGXYCGMeMOxbSom26hgEfq7IDlCiO+k+ZldSfZAtf6i+82gu7l
tnP12ol3d+i82HhlFyph1gfQN5ZIjAkQyIQTyPJIj55+hP/NAH3MoBeHl/oWiHKo
F3JmgRpJAKYYW2gSQaRCPRRA7DHkhnD4suYgKCU/PzAfvNu9iuvuDa8u+vkp+x+Q
iailIsfsAA9Ddgy7s+hFHtFCyIstyfZJzCTvSKbn+WRFYVCx8sdbiHjnaUZb0XYG
tjU4ZZYK1m1KWeFW3t+sCPfSGz5OCHxGqR3vXiirPgVEDLnV7a630AEdrIRhHEcg
kICaaYoYFNRlpYR7HeN+2w0qjn/Ntjf6jzSAjwibYYEv0vWputp4Pwqryx0rpb1E
Hh3ZHRq4VBDcjjXS4rOPembUn9qDrq5kSgGfVylODGNAMV373Yn1GqY0mUv/5kbS
NbL2Esx0nk8AeeSfceL4DqZ7mJcpY9xC0yOINih4KvTFh6RgiNK1nJvkWUcSIIpA
6x61vnsoP5jOvmAXQFgZaPtc95TbvQvcWAiPzmtjxAvvBajrK5yj2m45LOcHuXN0
6Ie8pcDcErj2I/sFKDzBGmFYCnug398WSlWe9X7nsMLiNB0BCjtfCnfE3Xahkkub
8kQ6PrNsuwkC0Ud+Cs1T5aqsXlMC2m5gQoahjOQiFCNLZzVvhw4t1hu3aDqTv5aT
YCfKIiQ2WTQ+gnkG/Mgm2zEr3xzpbHVNwxYSNHUmqC7vna7ihuVBMk/yC6dk2KsG
Q+6i6P7jAmUTWNfKbj3+WTbYgY8MyTUP9K2p9pJl3Kt5ZH05k8XCWUg8elLDA24U
n0Oysu50Scp/wTgKr48Dg3Xrib5xrQcNkeEAgO7V71wWKDNuQzDfJ9ndRP6oiI3C
8dlOzWJJZHoKjhivRFMiW2PQKybgTnVzsNFMC+nhmE2Q4kq1D5QJdRG0qvJ0TCrK
SagBfMi69DOPmVDjL0x/Tfx6igYzma8Ts0l81226DnqUfUYyjV4MmMKyJyq96iIl
ucHCZDgbh3Fpk1nWyTmOU+ZlvwBLv/6oMpig6FEO1kpivfqn1Smk/U0bPqXYwB4V
+aXbGOLF7J9kfyTsQxqk7ylrSiijg2ayFMUHZRdVMkXxDWXkQ0n7p8fNc4HWS+uO
2kZmaOw1MuztE2ViY2u8ISnE8y0jV/3uM2pUZ4heRtMrExOmXy9k+LOgrzkaRjXc
zaZ09oMwmzIkxcDkaeQarvpCab+MjXZs6XIA5ldKK8O4Yl+FdIbWPwUtexR79KN/
gpm82LZMHuHAlE16YooULZg47DweJVD5tD3y2MojrUUU3fcPrrgZRtlEgCYFsbPY
f9UxBcLnz1x21HUaxYsxQDFuaEb0jwMXNjjmgUgtnw+P+kv4eE9UfJoWLYa5dxao
9Lpsb3XiQVpcOIfKoe34N06IHQOGXjBgDRKm5u88lsdqP/dvn6+7B7EaRspavvsy
y4zfORRteTc7QHQ9Z6lwOAVFn/uyetdwCqkXpcEvd9M4vzKcPv82vpxFG2ErE8FF
CVwFlD0nzY7l+ms0O7C69qIapVKozrF4hxMqDTXPEj3cri9Xyf5lBqmcAGtiAHVA
5ktWCf4VKQDhUnR2vDrYzyqUNnyc394cEwoDRnAjAbHw4ECi29nOVGS5n+6JW7J0
Ub9c48QD3pf6uyXiuMxTPBor9wUvUhpJ73ZgXF+CQa4+3sEPdzRHt1jV1bJeh4Vf
BqseJk7YkrOTP6EZusB2ApU0yVubUOIIFktPsL7aeiEewl0um5q8XwGyOy+v+XMW
3dS5uSG0DWGUHSGYaiabWcKKpiALA2YqCkbKH9GHtq4T7pJzEX02/6i5C40psbu4
7AUVdBz59kKLQ/gMU42To6eWLc7y6Hiyz3TD0Pxx66OcxJa3gr5ZA0zM4UM7814R
PPFrMgcByIxEVu1BSHaAKJB5pmZvGmOo8h+twhmpR+baFbsS4G9GKJ9Lc686XBH1
rTsQvgGm9CeJYxY33Czq74u9s80xm6DtBJBAFarYlzYMdZPSK4niOKrIgYyo/4Ex
KpN1TS7pFIHL+FH7mYmEo7dtRH5nDzelbYhozBhqxTxk4Jru/XjtHhE4KKyvjIjX
QrUih14kqYfEMVYt9k6HXSo6he3RYAgZYuAGU/pYK7FGrPrb3bXgXFQXdJtLyuZb
YmqWjLEr0qjZSENop2W3lxAqeM2Rknq1z3Jt33nc/d6iCKTS4bLBZUs0HCUwr+Lz
JeuRdhJR48XprM/wFnpWQO6WqDTUD3OqUKf2CNq2TJTsdZOQwolHZvXQmy9ZYgXG
xkAIa/kuiTlzWMR0XraqYcKS5oriy3+1k2bDQ17vBLtH4yD4xF4RgNaPA2UN5kNx
JhybGDAZamHIoIAMGHDPni3Mh0aTM1kuQUpHTVAaVGC7FXW3JmRsy9pTltCVVD0k
0EmjDlqyOffJmqr018HjLtp2x5e5mSiyMsqbXgCBHr3b286qC/DjCS+DDVIyXKUt
AnoTsEIooTpn+MlUHgkmdW95WU6aDKX7kxmGdAE5nkmvMZimDqou6jxGPAAInD1s
+slNdABJFiazTHlJnyyeMReEKVCREgC8EFOFfIClL5ZOGAJn+rCnseE4VXVzOcRW
K2TPS5BSTgBZlGukxxW+GkM5pmI9Us3VIct0+r1Fu2Q/hIU1OqTP8p1+3i7qbhXJ
X1Tk6yRGOpVdRquvaixS/EUutQ0L24lwNcVxMDSaIgtoN+Lkb8SxOHEV1JubVpfA
iJi3lB8HpPXl2QKXNYOsnblJD+G3/hP3y6D6p0fyy9G9jqxz1582P5oKst2x+zT8
0P8oW7w0I7BXleOGeKZQiXWUNbz9s90SW8oYpeUUZnHztP6XBZrP32fUZ1e8ECx5
A2foO5ItL9QiQtnhJ+dJRQru9axkQKxVt9yMpgGlkOLI7OLZjY5+MW63pMFzEUB4
qTbXsyc8amE2i8SGBHHNWGc0gJnnV0mhHDCVSRkHMUKB8759EZpFrz9sa/K31HIx
b0luDjmh6lEGjrz3VBgo1x0PO+uikOsgp0H2sMyLshSX2O6w04Bndqmt/nJEAtuH
G3eyH5l6+2jkQeQk64noHOtqxpixSMNbPV31fxAWR5Dz3woDvKmyUH12guXTcQQ3
uEE/MBQaZftmeKvOAzAjKkOzCI4q4hNa+U/FAQGD0hHULyatyUWMk37TDI9nG+T+
1PqLbTrgmWm84hJNY5uK1/l5UOr5FbIPUFRg/YoKHQzwCuPtnKg+XijzWYNTaZz8
4uTovMcquebteQv1tCqgICAnsmjCtrUpSHTwgmJO9IFGpm72j/bwB8Up5u8ZTMHj
a8r5yj2uK3X4b01++W2t3SpcV3t+vtXqkiucBYtuu3VSqJ0CRIsgunUjZTOD5OTA
OWLMv7I+T2biwVR9vsuXsOp4YO4TjLFdCRj3WdJtfnpAD/TFq8tRYUDM3UfYS+BZ
7nUIP9ddwAW0L2TeVTiHEhPPUVc26HB26pWquyiJMoXIIezxFtyBCmsOKt6DJfPq
WJd166zAm/cUlTCM0ks322v3lZRX3AESP3ezl5aLEhYRobl4UvfmLHuweP2QpiMB
VRIAl+ELE65v606K+X4jLX0IxrOmwtkpQRJnGmXie/4cOnGj6wR7EVcJ7chsPZMI
xhlb3y6mQmNFswoO+pChBdfqMh0EKYhNpTDHKPmfMkJZkTZRgs5G820+ojvx+yl3
pt6cCfr9tjxQiL3RPfmQiZIM4qY161KDcWRNWbS3MN7Nt3+JQdByqVVWCYLDVJDg
/KTlapmXgbsKxvDl8WI6QDLww0soMfS/dy4emmuL9An/K3WJT1CrcOcsYYJTYU7U
I/LJylW70E6+AHtHTued5Be11rxa43LEJJNGJAbI0fFTleKdCXdD2Y6DMJHaVFlH
dj5rZ3/AwV7HCatSVLU/R/ZROJHeeoiCJZbPedf6Z9dEjomF/51p1IsIgdZb8o6t
vzZqlrgwHWHqV6fCGfJaqH1iZKVXYeFxw0ryaXY1TVejsW6GTcejVlFkHJTtddr3
Leu/y5Yys1j3zy8/RJjsOjoaJlcb0yV4fICh1FzH8VfvAPXABWPehelIAJxicwdi
nQcn0Rh8rmcVlQmjgAZ9iY+noGEjeoTHrRWhDv4ymAzREPhY0BaHfsBw5MU7gqYj
OHQAS+RnabhWZSUPWDk7g/QBCYzynccRKm/tHSTFOgfIoXTkbXH55BTk3PupUZn5
nCnswfxP9LYDLdcZ9Pacyps6IFMRvkzxx6XABV0Xq50Iy2GHmdYp82T6AOhlYoQV
8YfuyUGosinYLdVCkIuwJJ4cTZ4SsauVN/x9+sHGUn15t7ErooR/F8BFwjI8RQV1
kV9gyVBs/2iL29Bv1xiWP1mfIfNF/wqda97b35DEa56sYzPsLt5OzG+R5V6Ud0fK
f70EIG1xv7su92uY6tsYYT9f2flZr5bwQ9S7DIlbqeU0SWI0Z18lXkb+pqngMeGO
XwtnZ6stWA51oOyXqVG0JuYdc2sDT2/qLculpRrtiwr7qmNNIyx90yVhg8sSh7tW
RBNG4aSVdmaAVEwuRte6MLXCYxtQqRkwLlzMbfTjWv2n+d2gcw5oIIxDriE4j7uG
C0TLjAlpRPchaiPVyAjurbET4z0/Q4gMdS54hZPS3VbMTswEGfuz5nNofxEV0fDy
lFqDtSz8VbrwsOZaZA/Xdu41nlpu3UuyZLF6vwEXorBtyR/Iy9Bxb3H4O2MmigN9
TOp2gt6T0GT7BZDxJmuIeXhT1sE/2keUv5taF7qK6/qw8mnZj0/u5rv0rX6/p5LR
a8vXqBvUAEmEQtCFGnVNPPUlg1GbXCupKypDRAiO22v7BpF9m1IfNG5rhlMHteRI
t8CBjliIgRFO7yzH3OXCJEeZNkylPSbltPwJNHD13Mgawolz/R52M+fHKVaBkOi9
Xl52bR7zrXSk6ZKTnnQlbjXT4b8L9ru/2PSpxwV9qOc6KIpgdpGX1s0sm7yHLebX
dFqi/X92O5t/azcU8VGxAdJYZkhA7AwuKOYXF/SlXwmrI0Byn/Tr1FxuHjHytETq
ya/Oc/QplS2N1O/CrWqjmC93Jh9GP4dlkHktyJ+NZ/+DiKBbSr2c+8jLizTMnudn
oCsxkE1zLZzjgcMbt3h7hin0Ec31/7OKCZLrnwUqT7QQv8xJJOxteEPffQqGRxFt
ebjdGX+nuBPq0gKNQfgbErMepYYfywvzSs/ByTPOhMkeMMaM9b+r7DMoViJ0yzWH
u0FjglKmyFOU8RMuUWMpiTGSSOfokbIwPelpWXJ7AgdoNYKCbIXogl5YDwf8y0jP
ztK5XAFKNYxbqFcpMuhU+M/UAbLUAVRW1IfTk0+N3/ld1IFfHsdBoyNxOqV342Zu
cBrvXb3CpS1Jxn1Gy3XdYs0w1D/DoysDbAqrWkyz4nhvTH3ngbtpnRvLpHVBWVCp
aRNp2+hxuYWCEOY/CDZmJ8Ga3PmSrn8UtfH+lT0OnJfXtw41Il886fTbXDq/eF0g
+D+8VJqP8l3wkZrpTf5w9UbcJBiKqknxC481PISIZV/+vzaZ8ucyCkhR3J1MA1Nm
Qpo1w62PYLrBj3247Z63zLvvPXaZPDeHj+vVRvCvtCRnxccKfXFgzy3CAiYhZmGb
PyNmnI6TbQkMjzRtrD4ygzjNDQ+Zb2M5JpKfPFPjRjkaHA6xUUBeyRZy9jhXbO+S
xhb9XNVEJ/NV9EhwUaCGjJUDh/uiXcXnxIY1nUV5aIe0At54HgyLkBsT4hn6BHV6
LKrdCD/3+tU1ONQPsPE8BAGDoWp6m2qZouUnfcDKmhBy3j6VOwse/8lmtAfjYncZ
1TAhwY488JDVPEUZhb9RCk0m1coOmOn2dOmjlCgcNn9/xg++Z4aHGoIZiVfCyHiB
KVj3L6Gm0jRS6AT/EelB+i8l+6JRceAxd74YJxtqAkSo0zW8kqpXE/JLL6c2rnEj
qVUVtf2J6joPvH38hf0ujA69vnmD1sm4gN2Rgu4XHGNSCAFCtXiDS1zjj7gtuQuF
h/sZsYU4CO6YXTNLbAMqCZkxP9ar7NhAKXFmsG/k6PRBPZr2SCsLUXFPp+ijsxqn
9FMlj3W1yGcWkzv68Xzw+mo3OfrZXW0VbXecxqoaIdwwRLucZIC4iY4MOBAs7XoW
3LA0jUrlvxwBGmWP1bqxTzZ/bt1MDbsECD7eLpWAjbMuSCEp961ZOCupOFSEwRw4
dKEYWM5Ju+MuGfWv+YQ40yVdh4OXKV4+6NVTbfH0+QevGG6ToPRSMFu+eH+ZruoE
qLLrNRaklimdeh3TVA34aAu5UFb1fVog3t0vn4ud0Wrup8EQprd/jX+KOfT9KQWv
JQnf77GVhUy4e5i9yFKQj9sUZcECe9wKbwc/HxfPeBR8JIjXG41kM5gC2TucFu8C
7ZfEn55Kz1MCr5WUCaJPXAWdZL4ZsUEiZDV5TcBIOpCgC83pm+sQu9VYGpSzuAvL
OyNIIG/PpK/gMZc44jiPdGdqP7WXesQYf1pMUGu6gb0DwPBoQrxDiohbgQ6ILTLX
v8KYPWF31rq8gbsev8CFNv4dSPNmPrNNP2vjPdeea+7/APGibryt2+u94tt4mKF1
jYhhev6+gbBFWcwp+vPL0625hHwKHRmIg/nBBE6af9fNNgorc+1IJBlJbYKckJKw
U8gzoAA5IxWVOFyKYe3+5E80ljoBX3pLnc2QZjCy2w7l7q0AD+LdJVtAV30UjN8y
rArcwUbNpzsGZGOyYInUzjc8SMKMIoorOHTB4KDb1WDk0l0oCUmtauyZZudZOpCG
BxdeztViSV2JWg3QDtGswfF6ThFhMSxIp3J++/tviIfarCXJ+rrhRRYWaPCbzO0Z
+Nhyzvx76QaHtw1icIUW1YeuIhg/9curafJATTRoeJcpevBnM7Qi2iewqjnX7Ii6
kO6vcFkodtA8FXBttC7qXFMjkNv9qAj+6/gWOjg4snCOYbWbOM5Jwh+p3CsG08Rb
x1QMr1XMUiJ8Tgbot3eWit4C6xhC1JTj/GbM1LrsJZp4y+abQIrx5zxU5GQ9vZN8
KN0/BMI88/7i6Rj7moxirNCHYx5S/19Rt1zY0AeAQttpSMzuMXwLOUzxB6q+aEH5
QSsURGjB5jrgHR8R6/q/aFvu4BovOLJFncI7QNyWVzA7jaQZ1GeNE2Z/frabts2Z
9l2UQc8Qf/T6rd0SzCJWWRkhSHcwKuctcITliNEsDfbwHR3xTW7Dzfw0e4oG6uDd
eOHaLKZMPWOQcvz1dRnOZ2qImiIZDvyXFwt5ES6hmTV5oHJU4twsnbdqzEEm4t1Z
fY1yRIS64WM8snoDZaV9yjJZFiCUMttXZSm7dTKPc5FhreF4NzIba0F/8PNkuUqB
AyUOdPX0dWBDfgUGW1s7SZy++/N6Lqv9xIOa88qSVpomVL80o/vNWPqmIAuf0E3y
1gtBEXEPYdGxvHdnwNVrVmjc75PT46dN1pawJkJkTpQv0mq+EqqWDggqenDE9HyZ
88RsTmA6ocMeRw9aG1amxcIrZCrKBugnSNVbx7KtmIXPmL644tn7hPF8yJI1yNjt
bkED0KYbWKLbCLMcNq11y9oqb2oqOR/mNrFJAOklfrMHRMXpVcp1Nc+RezYZQcNN
v0SEO+YTN/057J2BYjmgh/2xQ+yPlVZO2KUiwOp8at5Fhwt34ebpOlTgCYOZSH5+
XNdQL8KJ2QM5WugTYzyzpy0+d5sVZq1jHvKwHXZ3NR+vxTNuS2Yo4muOwmz/Woi6
Q3oeKtDOTyIQOH9hu4lnS8k3x0jjMYHeJAAcDj9lFLhTNjL4yL+thzam0I8GnZ4m
RQlAYQYRQYmUcDgUg/ZmpSiI0GaZ52JoQw9tAulHvybI4pamK+zsD7YyDmYEk9hg
GpU8/lmAJY/7oDvjU1BOi9AFtoLIk/yGAj63TwuGvnJBBRWCFhnXios3+RLWXRga
DHKmoN6a1mNAfDxr00DjiqJKZW3eNOtPNcErnY9gMlo3UVsUa3dptE5ue+sGVRQ5
cz5O9Rxyi9/RiRhIoWjaIeMOk/1ahFqHJpi3B5WKn3wxVixp5Eliy2byFhPPdDrY
L2wWV2vjV18kPSz8U4sTrV6Naf53VD7b1ApcDcbxAobnX//X3bAJreg7Gc57WRgs
GSy+tf3HjMdEFAHdEPoaxnChEvG4etkC+k7plDy9Wb/JkrWQCdyM1GPUowPrb7fo
W6MT7P6ZRKhMohrD8cTyBCQa1YmaETXp8VXQCXbI+phtTb6/Zegvkez2loxDNRF3
dVOTeSJo9PJpGeLlBbKz61JByJeoPKPTIuyjW2KbGZLAT3mZk+/sjxryhR4P01oh
m85gWdevTK45PilSZ1vCyUQt4ni5UZY/5I4pDRGwz9XBwoiPT52auKUyL0jDr/ml
k8LC4mcBbxnTWvPCvixs1RXb1QnkW94YR5di8rS/OhfH3rU+PR7/02nfBRistgWg
JCB+8MxfSZ7EujmzCxVtP34kzrY7bWTULjaqquI9W3wOVvJhaCSESzataLn72/la
YC42Pnx3YTGgPq4vWS3qgpADqwbnzzMUJtokV6smhdqJZ5TbbE1oroTgaUMoKZk5
jwMw9W5siFnhavOa1FG62Moew7ITvQWTgjIi5P2wNpmPN91tpMJQYAYRCrYR7y7i
QSW1X9nrkHGXAm2r08XTJka9O6rcpHvrJAFEgnxI6dgF7ftMNX8NHkKxgQ6DFcPn
daXZtZw/2+QY28GBuw5LWYojbtp7B+90f3F22KByZB24RbRRziRjrdiCfM1WuA86
t8UZdWt1C8Nc6WmV4WNBVmd4nIu9WvpHJwcMr3Ji6tSJOS4+JRjxupoYMZypWIjG
WQChWhzM1Wej4dN9sqAhOD1MBPCVgFNZ/lghqJE70UT6V6ofwLJX4NC99ZsSOTeN
qm8a4vhxwIMPpcW5VHO/6D43RoIhdj+sP/UPrJ5TT2tKqyb3x6FsPYoxt1+WqYbO
mstvLWUD1Vp3RkZt7GCy9xUKaX5xJUi+Pr9LZui8GZ/iMzXfMR0zPBDWGJuZaovI
kRDMLtMJWTD6x4PTNeW6mjUpdewhyFuQH8PZ2YfDzo5FdIIGXfHsXH+2taupB6Ky
nbaUuW8e7ThHEOHhVWMjnb3Gv497Uxo6+lTu8exQZkMa8evkryLIzcPhh37sF1Nd
HB1pfASBrHp+R7liHawTIB2/90xSvWcxIYgiGiXmPsuNSnPT5r3xg3tQQFJQY+2R
EQ7oIzeUkZns50ui/LLwHbtsySWJ/ZNp8FbIukgA+Ypxoc5KwHJ22IpI2HRbM9Kw
Ax+5mr8SBUdlL5OlXTMHDWH2JJq80JOAytc3wwhSDWpUb4vF95LAWyac9jNPWWbx
0BAOKwb6wDFTGj5L8mcdRm370GNUiqVEuoDZ5z9BhTGqhg/RRPIkNdxJzOrdFukl
8r9HfsCz1SIA7+/1cPbI1fMuhZY9KI8EmNdCptBBZJqyHyh9yX9wFvU7epPfcj1U
zRc1dxvLtGH4oeS1QoIOgEECV2g+6+Qastmukbx3JHVr+YQY4qSlGKk7t0V3afBZ
++Zng0B/MfHFVJqNkoYj2Q5RgFZN/r1hS7G91dmHfgIsr6PrOq8S6VKUd5dwLJ57
ZTj6bf9s+UKZBN5i4uRKsTYVaPQ/9iqlmOSwoK304F6PTqSbB8PUCJ5BdrFbLBdt
tws3DmRECx9Lb9fZQJD20AGD++3dBiItt8bxMzkai8sgTP0UT+XaNmFP2tg7Vn4/
D1LgXqEdKsF4fGhkV6v8SBsa7jhrAXXj4aQD/IbEMRTaqKiJS45InPYxZ2f5i2wS
2IzFntQ7ktEGFXnxWel7vUjY87sp0w7Oo/DrSRBi2BIerDoMOMAe9MY+RCNrTdzk
14m5Lvmizm3aIUp1guR8egLnU0jXr+4noMBRv8ussqcDtwZaLI4Yj1DT5OORzBHo
mRLeQISzozWs1iy5RxpIxTKZvFzcLqsH1uS2owrq470FQOY2vQJRwvsW9oVbECCU
3dW5E2n4D2LTtYhKX+o0PENSAS3DQr2qQVHOgclZWJXjSZdF9ULB6pO0A44mOnJg
R5CGD8JjLryIrtoHCCH8+ga+1aEUcCg1whpC1uXIMyzFBHv4bi/IGk5DsBmsR2Nt
N/FT4GGyYrem2XYkMyazqlmQcqLUVnH4KeqGbO0nq+w1s3x2OmhFE2JbcIcxcpPL
maoC8CLJrUUvu45t37k6B0VhJtoAfGw/xmGOZ6cCG20M1GoRFgwPRUT/K4ZQuuMN
F8dfgBMDbgyCMu+DrQG5D3n7AH6WmbDpvePc1Astk3aR7YFEx8znTUC5abd7ttVf
6//fVAp12bxE0gTz2JkV8ojfY6uWrI3iL2IJAVGUgLn7KITC2lwDBBlFw8HZfvzL
EqLvbabZNl8ZrVF2LD+lzC/fsSkuC2maBfc7O46tpNJOF8EuQ7R1r5KUdqqIdOiZ
u3tDaE3OnsUyAmpH46wg1ddo1q1enfsN0iNfKDQnDKcAMG1MJfbbC46zcTNq0y8G
ibVXZdWqqRmMZavnsKkAgZ0u+g4lURktkucpQzYb/La+fvOjbDm2mdsn5nzJT/5M
GOnLftN+XhYlDEwYGP8csovkITc7A31DgLxc69qCTJew5fSiBuTtyfGlrm1EughY
Y/mAbrrKJIyj04LF5MGIUDiUEm8Y/8iyiTs7Y1NNLEYqtALIDuC8rG4YHNOTyZKB
i9J1eWQ6q/pP8kthByFkMLfDIc32npE22uyKc5IbfWuNNozta78gYkpFO/wKVpD2
FXUroH6dC47NmDy9bXh80KOEZJqhWWAYkwBmsBppfLDXo9xI+2NufQMY1xjSMWE1
4icduuZ37aoA/wQpjRC+oM+f394vkOw7VR0I+rLgv//AKeyfXZxVocsTCiTZVhYp
J5cA5mevXrLO9lCt3tQdQ5BLvEfQW6jzDJZ0QoIQmUEevGw/Oi/5Tldzc2YX0Nxl
MBC2nOKyuOdGH1RSFo4sffEfjN7rMabG01teyeUeFGMZuYMn5mvY2TZGJrGF7b1P
k59vhxUuNWA2Me0hoGY9oSlWFnXWb8uUxiHnmRF+OtYc66Y49x5kgORs2e5ttyvu
dt5Vq1AysmIM8B4s4/MMTY53Udy8yAm/c26mGaaoHQ9or/5fJDLHpe4XDOpc7rhz
weJBHV1f07PQ6QjviXq1Fy/I3KegPs+vKmU1fA3Jt2NEfCBlPMlqP3wgEsDSjfUQ
PuWetBC7Dw9wg2Lvm7pxjpeg9VWfXRK4NgJfg5kyJ+4xo6xcc+qSBCT2o7Lavmvt
gUjqunEAtrPS0YNKyAARZROhCCeHwxkCXkYUhn49rQYtoZLyY9ARLZPm+hZNVetv
rYL+eq6Yvkf99XCmXy6IQhP9dqyInouJmU36zI2ISsZ6Om2oM47Zu7VVgUlsmgCR
H0jQtEgen1jFw0R5OxqDEmHyCvXn8tdJFpW2UADxq+PRB+cHlD4mJ1TBaj8h61hF
zUIDF1TwX6ygKmouW/oBsqYbxND6B8zG0WKl5K0yc/DKzHaMZmx8jkKLtEbc2mG5
`protect end_protected