`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 27696 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eislOGByxcl/gRn8UziAa+H
mjgbsd36EQO5Ail/O6Xu+R+88VsHVstuDsLtmIbm0mEJbw0NbwNFUQIv8JcBY8vh
zVOLjFxuqm9RFggYxkRNNPKf6Jiy6mdNv0pV7eilaIi/nUNa9qD5umfdzH34XALv
aiKN9Ie1pyrqdmiqsp0mDXKXx4hObci39UhEO69ZwTXSCpN8lRyHlLlP5YWSPPwY
76+neQDxQlueA0CpWWxrzaShhl0U8dUj8ouoGQf+YnVEAZj/CGjhcWCpd47b8D7t
51DUQqS5h0UoQmtK4wv1stK1WGCMDeVUk3oqXiSCl8CgLWsUkO5Lwe5ht3XzsKxy
xcBODEzLV+2dKaAxJWus2sAGjSR5JeBTosN2MFYa1msSLVc0Laf7vYIsOuRjWi+E
bvdE4EoJQ5z2WGv1+ZQ/GcRbtvNp5JWfqNF4oUMmwXCLf7xiChrDl0Uo1BvHcz4D
QE3seRxVcIv7X6VmePm2jnGj2nUpTvOP5yDYbdn+QfnVDp3EeMPSELzFPG+N+ajA
Cw/IwEoWu+3DhRixWHkoh39e6D4ZkqneP5B0iqA6x80K4UHvuAVLSOzBCkTB0cA6
AWD29BBQc50BIJB0E93N5/orgw83Y+FEO0McOFDVAjkd2+qidrYxOHb0UaOgZ4dI
rErdsYFGILmMhdAQ7cVQboIIiyiZtYDkv/rUDoxk4hOPflmn82ger2EGFJuoImU0
O2ZMn96Pga9PEwfkkhjV5IcmOjMCVrtS4mRoI/lWOGLRNM/X7RbOb3u3mjOwtrFx
kDFh6/wonNIRLX2UsmV9xEzyM2jJBDHSoVluIQEQ4X5VePAgqtfEsi3AuHGxLStl
hM5eXNt+4jrfawxRnQbjabQlWtlyGD3KH2Zxocj58Zv6QXxBmi6/bM+RkF/OqfWH
o1bk3zJsuhEj89HYpgWC5N5PY0kOrt6ZWnrp/47UMBT1gmbGv6wygE33VzCbLsEO
UDwM0HHpHrOmshaIWTVs35DxQx9ZUCGlvblTp+RKxX8msoa27AY9iO5jlhUzgwno
YdwtFGzqHeoR9lCnp3crvYvl58kZG+N8h5RIpG6k0Ya/SwIEuLoA3sJmPKp2Zvez
tyDzpAH5NEHkT+L9Ppv7auq24JgcUJE1UufKROebgIkSe2cBWDK9PWy4hANc2hE6
8l8WSGDT6+JTlaf/mlkcUvUSj1foE/nklV3LWeRk0EhyOLXroyN6poMcsAhtvDkK
p3jpIU2foqhq3p7R9GanYAbDhtbXOW0oPL3bU4dSJjH49dyRONqjn+mYolNGKCFR
LcpPzdU7X6msDc24oub3/iKapdDf32OqaEMysO+DSEApnf5CYSDYu3AVlzfAQMlc
QjMkdQ7JsJ+jgPMQwEFoICet6V/WaGzXQxAU0aBrClUgg3lZ4NqARK5Y6ZX1ohzj
K8PBaROjxKEAEXxUuQXTc25wXKe+tdGsYvpp3IT5/Wq/kVXPImW13IZV1sP+fbOp
y+eSkFRa5k0miZ3EzKGjxlVzfPgo+jao1ldb/zGKQApVmLfzUbqHiBIF9DVGI7BS
RLF7wCaeJn6wr01g1066Qrenh4Z7vvXsdAzxMeieDwJ1os8hqR/dnWuAjFlrjDza
/wuSz7OVy2oHXRkAsEwZn5fv7huZaATBYZMlC3dn6ThGhG4ds7icnl2Sgt+8QyVf
ZhGlQ2KWMLF+K/gAdd8URrw7BPuu0cMwq2fbhEwG0B7dMltR2vjmdWrY7uIWqpgU
E1oki9UiVaePNWHN/mT7D7D9c6uey7x3epa8g0pe102H+LsKVDOSCu6aNWuH+O7w
4K//pTHxyVNe+h98AMly9dnveCAOaaI1tePwasyU83iC0lMnaV2GbvhqZ7gURGhN
LR65mcOxiebq6cIs10OO1SQXMpsADclDzI62wUn6LJ9AHTZWy31VvhsG7AE36HOw
lm3F9hE5jAotANkfzaKuXBDeURBd4wqEeblYTdoRguio8BGwcVngrHfDwIZ/IvG1
hFJMIIPs3yZIL+zuaCbycpTBBRdx/JiIy+z8CzZYYO2dd2JcgbhiRBYtgUklBhqk
woGFqWr+eph/M7GQj2PKfBjN0aOuagb+bVXuU9IjcVBOechrkVFJDRIltrSCbi+J
7gFzygUWlDYgkVwgnxpHq1khjItUSNl/noYUeyAP2MTAQDZIfIzJR4Gj6Ni5iGpT
Y/Ki+Lb8cLCIQq1vlrh/CJBUt4U/t2dbS21pM7xTe8EOfp3Xcm9qHUszplr6KCcH
Kh+s3pAoYiQRfS7M54cbbq0dL1q+L2mOMdzwP/eGhNmYgeAko5I8t8meJ+1PjWiU
XFLwGakC84PHKxgMApCGkGk5rGAGT5hjmLbQudWHQ2yfleJENAhQ35hJ9tjmsehT
0WYJuuG+llYIZq547eiyyHfeIlNmhQPOOEOREsyi0V1FL8uc4MJANTDhwbU0y20+
PAxlkjPHyOpHgO9IY8DuuMwLrZbSfIdu26JENYNZ9btUCM/0gvxNB8SUEfDiyu41
Eg4t5cZGLvAK3IP1i28hct00Ck1VORnWJrnX8/dHwfcyDQpd2BfYw2+jUp48K5u6
cm7lI/0Dwg8bLwJo1VZbMRfU3ABHJGkPlVlaWKv3McCjJa3B2UsHqYAKHdbKajUE
piof2dudjNac3w1lkEQq5WedoeaFVPplQg9sDP256KZn9iA+TKGucZAih6CT4ljc
bLBKKutc2DMce+vzb+wilehTufL42RSpOCWmaOrVZh9HksVugU3df6xwrdxfV9FC
a26ZvJdLiBg2G7GpiT3Dt3L9DWbmGA2hCnwCTYjR8xokMvIyPvGF7P1vIWvZWdvp
FhWzmnRK8TNK0n7PpxBXZVvKC2PlsLLzPcqA1vYz1riWBV72Kv4g/mi0wh4xe/HU
zBFFYe1HqRm4k1KjsUR1bvN6eJ4H2ig1aFCgyZetCi3l6X1c71w+ux2h8sHTvHpm
PIMs0JBt+GeZYOorBMvD1r5SIVb1MSd0fE9YDChGlSZrjbl1U4XMTccNilgCzT8C
mik58g8M5EX7dcaa7YZN6vnX0L5AScc8u/HCHzbD+8D8R+zWIelIq36AYoZ/YHF7
vsnIddATW47AgZ/eWeqGHlnH/HxbPazbKV+SIl4Ww/8CQeiT+t8sJ/qQgPYposUB
DEM0F3xa9SmfvizSbkzOtd/wizJ7AyMHm5792dsg3xujlDnlfQfxnp9PfWW+oSLr
At6zXkVxjNWC/aKeu7UPHsGa94Nv4rKxXpez7G7aadJR7FKUUh9S25vgSOVJuZyh
50B1YsmwNfFx7rbeTTjYBxP2Xk/io5gsFjtgdyNI4x9BoHsMIKmLIsvlH2znvXZT
swRWoyXk2ZRXKEO8C/MnNtxXcO4sqtI47VdfCfP12LidP2t+k2fouC+h9IbKi8E7
Qnx7VGd7XjhFVv2z0Gks8pgeGUBCoBOYFAaRLffvzC4aWb0ggcb9y4jAOr4WUwK7
3M5HFiP/d1lf9lvDd+dI+i2b05Ee1EjkkeSuSaGCDWxY9qt5EEJEjTLcKsBEVW8r
mMEwNyaxajk4S9utPomVgoGWxQrOJp+m4cC+bhtK28H6sU2OTA0BMefBqspqKrPG
sguVmbhq4Ai5AThCMJe7yOcjxaqYhHO13qe+DHoApCX896jo3U+lfz4x3JsvXdG+
PT15/x6XbycbStTZeEk1GSz0Rbf7LVey/jZ9Kpl/AojxJnKMTkT7sKAfMV2pLnDC
QkH31KCJBmm+PWSoz1DExTnRFXm1La+3EmlLamd358VFpsMAlAJu9oRcXE/9X+1O
HcE36iUD0IoTalE8uFRArRLhTaiE+T9I2SXSVBaAXYSWrxvOq9mkN8u/igWyy/aA
P+zSwQXCOyoWuxQvZ+OMeocwCsAEQG4Ski3ZJwjw23gYp64xiu/JgwpTZbWCGLHK
4p+J6slYm5MAHJrEogB2zbTBd7/Mq3V4Nj0EGUaexX0PCzCuV7m3Rpykxtc2DFw0
o4MfZ7Z6EJ4LFHvlHoV/itQiX/WU7xBp1N8UTh7wJANbHQDEHnKMQR6ZjTNwQfIf
v9ogBSEcy8OqPHfVk5BKdjJGeQCZrOkeVaCnlSkrdFlqfrdhJF8fmZse2oV4I5Ai
BmjWNT+w2aSYfhqF4T12EDH6XM1+3ncZNIIbOaDCCQs0rzshXkU169bG27tr/SlA
Dl9bRNbBra1FoR5fp01fc/hwNt+T8PtbWfq8VqRCz4AgAbSPDPB3AzJkStg6uger
eEXT/artjKsI4buNOyMboKYUtGadGxV17vf9KfNyMhsWwMRPjAXyHQybn73KOfU6
3iMnqFMEJ9vhceZl+ni0NdbgJG8lFBYEgfj8W9W49IPV4rJkbcncEyLJVVXx4SbR
iyB/ngu9yUcsS5YOsJWo2rgyf/LYvz+OU6asdu+0FPGq1kHkqES6I1Xxa8bPmHVY
sj+ctr8rP/P3QSSOXe1bXBl3T1f+fnFSgJfRbuh+QeSb/A5/N6Lw4Ofjy2faTg9n
UAeKfgCfgNITJssND62IIAdiKXVdGCOII/kv2Pht4rcteInMjrT8Y9FVUJhgO8qZ
8LAZod1cvpBKDqAr5DoV94dXsdR1IQR1TjpGxmKZFf0KrIhKAyFMD1hm/BYIENaI
PaqZ6n2ljx8TvEvh3/+6qlaPtaj4rvbMKoc/RYtr/31Heih2D+cksjWHRYuXsvRJ
aXgKhGfp0ct7MtohXYZzTMoeFmlFCNg0KMjr60S/7qSHFcjpfZksQUG4vDGhF7OJ
YtpeHfBJ/u90H1CuFdWvmX/vmKHEKEZ5qNGXyBaZ7Q1kZif+L0R9zX/ncouZWVKz
4gobWpskOrGtQOIPp9AG54cD96vnOMOBkduUxtY+Mw2iKhAZf0OZ+pFeA/sYACaj
Bm82obl+mcb/Wsxilowp0T4vBZoGL3jAiDofBE3ujfumfRATimIfNSiPgWXDUQZ4
FydujVLIFubH6h4VrbAC4KJdfM38aUyTGGSPSX/nXD36oPLrKXiPpWhhUnfuJCjS
ksqDrXY3loOwk0W/jLCE9KdrXrIBsO5IQlBBwFaZsUyWAhTxQhOBvWckZx4NqKmp
vyx08YkfJ4iixCwTQLBx8d3QxuCmp435GiATCyI2LDK+0VaJZEajt+xMkj64OYdJ
m5LWltGpXe6Qph6qDGxWoeOlAxoLRVy6A+ibJOfOATrRktXMqDp5Q55+Sg862Hv7
rFt71UC6pG0m1NMTw46AL9wegftzbRhdaj2AHRKXpFmJBvJamWwwWsvR71VX60oy
2Q4O5B34Fhwo12WykY9k2J5LzfVixbpGlUekgB8xVaaGT9+TfIfUMzosRULApvTo
Y6p2MUxxnh3XmUnNJ96kaSVf7iQc+VzBpl6b1YtTknS9en0aKRBK4p7oXHKaifUP
N22VhDLndW5kfXAPwlP5PTeedgqvemw6SfgZnaqf0CYRpsaubYZkGdASgbHsKkUl
JytK85aZag09RPwPxEbAain2HGPTQi8qr8MLBaqxKZvLCZySiQ1M/1jM7MXllkMz
Ht0IMlFDl5HnEBubjPql9RKqH+H9Y+PdWS+TrxF2hKGjW2Yyo9eJ9v3VvlGTW5By
H977nmGagx8Bbm/Y87MqNp68bKW4C18A/g0VH2EQAH+E5Z2zQlw3VGVMYH62DQ1e
+UgH6m8kvn5t9dtwoK6hfJcp+dEXrt3YcyNlr3Kyh0viEv4qnCb+JpQYPhCRfZEJ
JtJufw/UPZWRFWsg0gsFoR8av4o96eisqCxQXiaf9mDnGlb/m8S8uQG84GG28MqI
DIF/+bQhscTwbae9wvJxA8jhhhsIXdYDoRXc9l5aAVn/Wo05ghkEsyBmYyQu6nPf
TH8j79fo/Vn794KWRIimgcWnbCVURyG6lDZjkIPHL7D1UXN+lXoB5qJ4IpT5++NU
Bg0c47QlIw2ThG1yo/KOpfDcCm7jQOPsgIFQAVl7qsR17jHc/wNQ+lcKyjHVh3Se
BPmxCJyxyOMPS35NPldCBkXeOLm2cIO26fuEduuNs2Ft4To/GSTljX7aDBYHmMgt
jiNglN2Pxxgc/aAjN+rHd5ipMoH+aHhwe8EYXJACer+puRYqQyTz36jcykpr2fUm
sBWXVnq379U8dg6mhu2LnfTrraIRSS2vvqWtC9UgOBfz+g3gn/ZzYKsqSWNAGxNR
t0R9naD1a2xJpXImYelI45FPTHXlgomm8/5QBec8ObXFmdQbYE25/kCaUEgyTjzP
gYCXZrVgN+DuIO2URw73fBjTyM8Cuqpi/cx+bc7L7P3L6F0Dzr+0AUExEIRigAca
A6hV1hGHI8UMIK4RBLkdAQOcexbo8fORCM1+hmCKe0Eb/rMB5ebt3Xy8UbadSl9/
w2jXuRcy9AXnWUUaN1xzuTNfWH5CZOfzv9kVQAW4Tqk2eVr+KdgU8fJ3/sDZ3ONf
LUSOjQdX+NbJ1VNX/eBuw2P5qFpymKKT8HWE+Qwzm0/QmD/Lfo1QzNL620k6+Xlg
1qq/WQbJpfPBGcbMXu4IBkDf3RZvNSurqFCbGjzEcvSrFyRC/G4P86YaR8P1wPEU
jLIonaoYzE3V6MXVaFU0k8CY4kn0dvoFbDJc+u5tf/fxXNEoqrO+217GtwUx6obl
Ikyq62I1lYCzyeZRvD2Ks0RyMUUbWkum9Jyf1PMVD9Sdk/X6qCPG9RnFQWCSejXz
lpvrMLRijayQBbuSw3umK+CLlMTeHUCeVrScVBRO2lrCF1Oi5yrDM9Cru3SFCxzr
33dsej+o45TbyqoKR/hL1t7Vewd8ZNRKHLX9/lcK+yXzYZ9/ypkbhTZDDsTKu3ni
jWfPPogRcyCxpWfMtTe51bbjdFekVUW8V46B7zWvxjH6UCDwiW6Tqha0x/tIrmRx
27zfB3JV6GdpcoN5eIg50qLUfVJNZZ4swRvvC+UsF21PpK3Ydk9hO9/eVazXe5ol
/kJZZMZV5W5q2f70wd3tkypbTRmyxCk/MrRsgNB3t494gtEI9fS7vhtUglNhakqu
bA5JowNoEYjtlr7hHivNzI2WrDwaZmEjG+NOVhTaAV1NOpQW3z4hQN6kUn4UK9+Q
rgbqE41nkE8WuUlzBV4f4aHsffgI5HZ6hWPyFZbP2il2Y6ikXuTIuEnXjrTkUun0
1c/pRHnggjFCBUzha4yj8qKZeo5RQoHs4+yxtvNthpYcahCgDJ0ysHoqS4WIMtqF
B6JY4JrqwL4B5BJ7d0Tv+rBLEFA8HfwXWzBUeSiULyd2VlVHyjfDUCjverW5s9Po
a+MD48+FbxLS8YiYwV+Lm5VeRh2OA1h0J3dH27w0iq9rcJB+UhrTJeqzULOTTXkN
BzcmJEHuIZnSwpss9nkAugtE/IMFx85ZHN+baMfu++rmiUFPUzq6oVwf0CS1iiJ4
KK/sNi5dVYtCTnU+A7+U1SrgBGRpR9sKk7WswyeCR9z3k36ALobY/Cmq6ZTvlQkQ
eivdcpYNrZpaqGfswQmVoR+vdrIVuN/F4Qd0MXKI3pkSyO25NKuUXJFxe2Bkw1gl
dMPys8hv2gZinDK6I/PsHgNeuEL9YCdBLl+etRWHyih478V+FhzWkttGrvRS3pbP
jZsMqaO6lrVcmQ8Gn86gvGoifZZu4gpmylsUE8GPHS5LxolsIt6yp024Ry4BKfJa
M7hPVx8+exMbqSWUm35GmaqxuLKro2Crbp1oC0uAbBhGyY7fbCV//ebaXb5+LbIu
UmQZu51WdCYR67Cw/iZE3aFpfgAuzBPcL3HQo2lQr74F3CAu1OqP+junD3KIo6UG
t02tPPowa6948hWNKT6PpJTRYJAeuofiByggKONHyOznEPZM6mfgitQDW5cXHQlA
LpvQx52BsD7CTmpPKtph9RPJGTxFtd+EouaOvhLNP+Jyi8FxP4UCnXbYBGm9KMS8
OIncDP4Mwi1FMsowLLsM5Rm4tdczXIobCcggAKQ2W0oacxcs7jkEKl1pnxkt6aeI
YZz6bPxkqgBbzyIwp4MUbIAeQSqtKwcfNlJT3+LEaf32rMagk4iXvgAegyDmOP1i
MRvNTZ0Q9JZmAJl/+HYFdo9MXL7rY0Ls1PQq8XO4TFMdSHde/T9WYV+eDgBSXocf
JoeSBGjhzAjEkmOBRPucIbw2iRsqqbmHewpVdy4MpV0PUmN62HNiQn9lRqvKcSN0
CZBcHwigwPgMfm0U8VlqoD6BIjbt/wU8IqcIjylUkjTeOk6h7ifAqIU5WXooxk41
5n6IOxuOqSOSYaLJJR6ga7XlcUaJNxAe8JkcAYha/+64vAV5Day4nSKDlgkVlfJ7
htyE+MZrelbJ3fa6xZrJ1Ng1tfWrrkjogAJ8W3h7QcHXyix3lE1Ag1k2v6a9VyNa
+6FStNkLAN2yY5Pjm7AYSP3Z5E3qykgYPuI/xYntbTxTQHPPhO4tvB3m0Lm8RHhj
nYPWQRW6yATgXWF03Vw2BcYcYERUnnmU3rU4IwvPjTzZ+kOdA1uBZR59ecY9np2+
4D//xdZeW/2jwa/2DY3ltymZyaJTvMiehZANgXBWNO9tURL+BtFxyzetrdbhZ5P+
LI9F8gC0oyEpkAeioPhuSTFP8VlFTt393BJEQU0uWBtTVXRCQS/rtSsHcLWv2VTq
8p8mjk1LguRw7ZDZjy/t2xqHyBCIVCR6uIV5Ty5Qx92F5o8dyweRSCNzg6FxRBoq
/hmfgxM0tClqitsmxBrBl7cSLSsUyKbWPU8bG6jqMF7+JJhfgdwPQNj9ntVBUc8u
kBcIWsjWs168YUzcRjYzSxBZbZj/LYoc8seoby2v4FKhWV89Sbc+1NP4HyX0SRto
TnHeIeVNyTomybt4sMqgamrc026vVF9GyOcKB29KyJAAYh8/hqprj0eJbxb0ahlv
gv/0JGskZEXKeok/sT0ZLue+uoeX3S04zOJRFE4MlpKj6InoUqcvXXDpObR4vc1U
JWLj9JYFRbru7exN95FHQTKS6Hh0miDJYWIiTrchmGN6BzWaDnyaCM9+e/GwVvqf
jcO/fGc3hcr6C+HRORLyWYTP6RdL+LhDKejLUaFZLgWC2+IPxwbDncsP+qcp/qQr
H0QtCi4Lbsz8x6IWBdgFz2vseMrHgvXbIHA0eVTVQdlUmxCJv8MtWJYGRwXcYO+Y
axuXC951+RLH0Eg6wPLHOLTXKvaI48VrPrPP4sn9Nvr4X5cIpKefBduGFe32hVSb
CxeybD9rY4wslaUapClSipbvFxOJbELnUTHWNrvqENHE5DeVefu6T1UoeyeH6iPX
YCOXq5py2F8GZ6etZQcoSx0OazkvQ2nztmrKjiQL0l2lDKuM6EfRsWRhu0eRxEpy
Ensy6kz8yJctfLMm5Kj+a7tr15NH0/++gnhXlvL2Q05VErT+cH3kNHrnURQVqN+6
gTqjNseQsSqzGV27ElQ3WgKarurSYJrgycr2cpNLjc//J6g42An6e+KggjzwPdoG
UDDfBXGfhjExuUvEioM0cpAioJIF0DMtTBXjrIhQxJaWbokCSkrl2jn36RPF/8C5
giANGqEwoZLSpsiNUO8JndlhsfnpUrHsu2IL/cFbl58r+hyiUrkRXh34DBqoPG65
Ap9L8ZpHZG17Cr4v/YljxSvV2zH4YQXMfVih816SVXphgv0k0IcUlrHxrrwma87j
EYtovnGAWXsRbnDEPCFWEackHEsO3Baa66O/Teytygj2LUs1t8KOY5OgUJIYYKCA
ew3qfPlejVLKELXR6c14qWTwBa7fHsZ6WtNUHDquADes8teWSRlfo3EGyKAT3vPA
OF88oKSu9cOEhj8n3J2DkXaW0kxvzMN4kcoKZWJvCXDPzHA7t5TuHG9EVufKwsu1
8te99XRWRsF8f4AK0jmT818oQCycB+EBq78EBrKHzLv+Fkit+c2l8owRtVh33Eb4
9pbn03GpbSPFza9zqV4BX/R8TqfHntcGWLy0pHe9yVADrK4OQ8BwFLERCdm+vwU+
8DZisACeRmU4T7dBs2aQG4ke9HU5OhuuBkxdImW26Y/e2qeEwd3vmYyq5i0CQITV
hGWmmM3smRPwBngyuARMhxR9ncigJp5T6fvS1xPv95NJHdW/vA0snoTQ/fkloVMi
3SBZ1f77+yXbpPgrF1tLMDfyN13bCuo5iQ075gmwhJ10midkU23akgYTreEALNFH
yRjA530XLonwIm/JLu34dToipVV50LhWvbly5GEnE2eudYCCJXX0HfHHfRzbSNZJ
XxhY9YWxwOGb96dINnZKCXdsLNBs5elpFp6U+fShsWMN092FX2hK7mO80B+5dGKV
Euqx24q891QQj9ueheNd7z7spopr+3LGDRdg9DnzUZCsHKueeXMC5rjRKox6En6T
PG0ufQaPhlfWbbBJMUpw1LUpJMNpnfc/w4NgfV5Bn67cr9wcgz6+0u94nkR3d8D8
5bo2HSOz3FhWJMFC1tTSWkKGAZAyn5aiZ09ppI+87/AwhaUSThvqkUK65qKVOd/C
KDZ7yxLJ6dZs7jIvu+Up1J3fKUKGfRkRFJ1h0+MGlaLPwj2xby2XPS7H2a303e4z
1ahfxQysBGChkTmLDN80iF4/9MgM+vWEhADoxplFdnvcAQLVZi4vTjd5+iugNBCn
vONGcVlWyQJbv05G4Tcbys9nuxnR913ZYjnMW18g56NwYNRl54vC9A6fR68wUH5x
2zheP4C9FZUTrD3EVlujBLTHQTHIZNENvJ1Hr62hZ/prhVkSzJz3w2nHHnIL7ax1
2ltWUFc8lB+vW67YdY5rroJZATXtRDuNrNWYZmae3rCeBGzAg7wTWum3s9TGn9Mv
DvOFiNFwloM0TTAMwDWBsSHyD9U1oTF8hD3wkmzprYwl8sgjdtkfBbRDVJwxLfom
PHl9I6t/csvX2G0/IpE+R+XXrIgD6Zsr/ZnYZnBRrrsOJ1nz2TVjM5E4ef2+AxUk
+UW6uenHEUqCactlxds2BqR9E6/PUBuR+ILMp3cOIh7oBYuAqOx3ToXRjWLQefbr
rq1dBKRhjD/ChveLu96nOa3WlxYjuZHZSP/AhpuxjuaVPWmDgjvMElek5jZzOsg8
uXAPfe6iGthfQTvgSY94gdmfEB3UvZuZfBVb3gwEEqBPXxdjp1AP5dC1zCT9sh65
ALT06tL6m0gw1SdUkJ3CYYBK1zQrAI/rwViCmcgRbe9dwUvmsIfijhvlGRg4ohOL
Dgz+ADf8923o997WXm5UYxb3e8pA2Vr9yOSi1lsghH68Z8Wxq23TI7MO4djWkq0/
pb4dnO0ZDz5vSyAbLo7vbAhXtBTwu/rpgkHnBDX/EYO4Wr7BbibBFbpJyDyrrRGy
kXHvhvpoZ+RWTx8nvh9CBi9Uz2RdArX3kst3JuvFesn/VImb1dywdOlJ+JXzritc
2NcvJ0Bw/69FusBXbjsY0p4p6GvaHJwaWFFAjmVqF9txrI0aBvUOCHvhbRlefYui
FLE4VWtsgUWwEW7tRzAy+tXSeWyjK+S4yN6zkNC1ABJaolpHR+PgbdMEERK/oN4o
EoVjg6PpabWHododCTGeTPPZE8khlawGoW4GPaHhIad317f27L5Fnccqf/O3NmYH
9yt0DHNDkxc2cCIodxOrW4D/4EY7xu9zfhggshba0+hcMgzwCJeyhXf1Qhk02T7j
JuCeSEhzpviSWRu9DFaN2b7QAtDVSTDXdpwzLVMMt2RxNJXvYiZtwZ993ENoduJh
DtHTha2G1l7z5yQDbhqnxNRSudyTQ4PDuALi6Cx63peO1c0V9IDe3LnlqqeqeGGp
Y54Hxe5sz744hKuJBtOJINHZIg/ST2hAuhU44KQIwlU2ZI7oTUf0/LoI9htvo/n4
ccJiJIyy1JWlHwHbNGoJgnqYzMjie8zh0S9SFPCrs18KHnAMUt4Fv4tNyE3wZbOS
ak3wlIcwcyk5jXMWpNYJLlK00jGVD2KeCopj8gllL2k92cFvnDUlwDkf17CIHo48
sPenioOfdOtOtdm7dVt7Kn0tzWzZEjTkKLc4JRa4ctloOu2zg91KNXvbj9rmb0JH
TtxqqSp52b7he8VSvcRbEtKRfLb9tsrWY4Y27GZ1ar4LY6ACmFSW3kNKtMRmu4D5
L0hS1tG7whBvrcXua9LeGTnJJmy5ugU3hpl11QiMXSb03bgoSxgdGxj4EDyLMlWk
3glJ9SIDfNB5WQ0WDA5T5bw1W5If7crhjW7FYoC7gZVcO8b58t1UM9j+zdDjKaIG
/EuTZtDncx8vwaEvYphwLwAgpJRfpDCzPLLPux+aV4dBcGYTK5+66yatRYb8jvye
N0ZWNkyO9EoAAoJC8dz8Kuf8jgFeq+brXTjt0UmYnnQs1KzOY3gDZ8v0KXO3dIhC
sJZUZqcDZaTVfh0vHKfmwArpLuuPEjMfb0hr9Wl3S5C0q5k5ltI+LQE/CmlKfRAO
G9Fin1d/SglsUmIP3pdZOXPAEmHXffoDsm68R4ZNmmpCXTnA0CAILqVvhEe/Szeq
XF7EC6HmaHBjppjlEQdoa7kEEewOU1+8/vn41lh0WFpkrTdTk11jaDt8F8wHYQ2z
X6ZReZIiB3S2C6CTaVDzbmI0v+iiof+WbHlJ7/ud306nwdduVBm1l1rcFXTgYbVO
PzCuqKpEKExr7mESpczX2WGTrLp7ATiXG+19Gv9TXTx+tAncFzaItl9JdqNJBawQ
Gp43qXj5h8gSEGSpfKDHcEk5nGCQ3bR/NhEfpviIRrub9/TpDh2Whr70PfSetEXi
OBMllnQViIuVPid4i3sSlxifjNrTSbkJ3SLuxsJ0alHEsANKmF71QSJ1Wx6WDA/h
uz7dg8YY7YENPOMRPb8MyJQXqvpxwPWheEDqT4HiQItiikNjCtTM+0pZr+96zxOT
cl04Nup1C4eJaBla/3NHs85ZA/6X9GpLt9kXdEIyWCLeEZHkb1jRWnSxG+XK2FrP
VgnejTYZTiofm3ySx2gLO0SKOllrlhDlYTIyeMElr1kvJeFbshBr5KXpRgDkjlWH
jTXM42+UGRIrY2OnU0y1IkpHT0aVICU0Fn+qq8AeJ97cXWWKPT4uZ6vGFKCEMFBa
QeAmtkz2gw5dK+vO1ABLxUFUxHA7ZFk9eTXxeyHqKaFT65XAZRn+jjt78hl5IKje
XASp0NZS3DvomsdHdtkqAp2a54Wvb4oT1pvwjeG7Kbqm9Qm3RFz1gFsxnPr41Oeq
g0p3S/sEPLb8rMWl/ivzV8qa2c6fDQe1C3xjQ5Bial5SUtfSZreJfrbAgBDxDFYo
rI64eDbyLb7IMOMa5rxhL8YErF5KGxk3OS6uPGZDANsZ/BbpwQaOHzHNxVm+dDeL
Rj6V5Qc4xlINXoIzqPV1yES3cmF2OsBPuMkDBMdZITGIpsKONzSVz565XPqgzmRO
TcV26Nj3HEobchzrpKtK4Ze7S/35GTd9AWPjGu7sxad2SiMFR0RVqZ2E9MhUogGy
JSVoPVjU9fPv6Gr+qLlsX1koPiqqy3bx7D000bx00muA0HM1v0VyaaJuCqIE+YbS
dJeHF1SU11inRSNbbVXP+vq6cvhwvyEIsLVxIwgq7o1KzsW+/NoiJ//5pv8iHm8o
RcqCfnfJKXhj+Tm1VcjfIjSEo0PtsGQSdaSKBdvbnwlqRl/tZMLyXdxSX3VrrtIN
c0/eJjkbNV2GuETLbDu+8Xt0oCC8WGP/JEKzP5c5M9Mq/Ivg4SCr5DaTWMeDjXxk
LeWa3r5MZWiz6m5cIhLuCRZOGpkX65LR892iLqC3C+BbPDo3deTOApiTKNhx18/H
akFmuInWv/Ghq2gKAEV5uJpsJIK+Jy3qWLj05FT/D0Labu7wjdhdx6NNoJYv4RtJ
sqgCE7ait96OFjE0EIr04YR3nAFDFPIPiZswn2dudDFJA3T0WJOuoexTyJbfg49I
TTEBKhygDBhF1Z4Nu4RfSkM/Ycf/n8ykYsL0cP9svEfwaYJbivGpVx801bzH2ilb
DR0otrigJ19nEpdoKia4QIF1DnV7NgzJn7J6RZsOEBzVUI8GtelGc/D4isXI2Nro
tBzv6wLebMFnl6NmBH/Gr1vDHJBMsxa2YXdrsl/5Y2ZA8z2sKIHjZhq6SUoE1UVu
Le1G1E8W1zXFCo0fDhmeLFuFHb3X4xVrOgVimmzb0bGaSAS/7FYvU4HNbbYBhG5G
VoHib3js3YiQc22cUpY1kLeuJD5hRY5FHfKC46xGpMgpzVjpp5Xke3iVpQlXBnFv
1sWTbP4cISMjn0vgMuHWFQddfyEB5zlfKPxXkyW/1K4qgWTLdYrmHiyLQVlVrpdV
pUiUyUdGV6fJ/gYqIsAXz/Nabp2mgPIvVqo58Yej2Uw229v5G6lKdiw4+Vj+8yMz
2KF5lLnVt+xp0EjH3jyjWzFaIS5E5ecFFEUCE6Qom6PkyBF8s1UkZV+26G7acoKa
HAQxsMGK1lCIfY6/3xyH0GIwiaZTQEvooM/BRHMK3HqqGi0RQv3ORgBTcLrrL///
6iqKZ9nuUQFIHWj2PbYVfszKHg2IvSzkdYGIwI6+1ASvYgS+n1o+Yy340leoakSh
syqX0hkrVcjaD+D+D7BWORCDyxx6wQcSQMGaoim7E6CyzIFTVyKDNbmZ8PQl1p8n
Wx3B6Sc0U+ZUWgTU0jmZ3umxanfdeAG/zYLrAkwbM6DMS0itx85OkuBIZtEWHQ7R
iyz7GK+PDi5riI3PRQoFcYe6LcovfLKPRZdxkz+6WpCUZX4ie3nvRhAAWxy6RF+1
BnTdjXL9UscfqVvUzPR4QILcKVvLbxKMkbfWRu6Vc4hpq6LXkZbYbGXHBakD/Jnh
BZxMQFdJM8LWCqRFqjMZaGBvZVSI2eC1dSx6D7Mh6TJDR9xiBUpDUFWxvnBldG+n
NITaxRUUcC4RROcCeXlusx0G/ZboYSc1+6r1YRQsccoo9CLIrHUpTwPzKCOfK8Z6
TW7pS6iAC/SPF8XCfBki+KyYC20nFW6YPYEn2EcvXFNj3ErLl9s8RyGUyPnH/R6V
t7d9ExdJDyq6Ob1MSt6vV7/oeg/rsdv5yAD8uI0W+2xMnB8CsDcI/tG61Y6XF9tL
llueoBLRL/qu9DF95Pj4SlMsDH4XW4FxZzq9MAGPJFTD+NV2BRo9RnOcLO7uY0FU
Wdv+I6ApaZtPP8n7wwVTQAroJGMPltQcT2E6hRleswTjJyCmHjELGgL874N9dwgQ
kBtwUQAUEu7daUYd6y1xFCaZ/OUiux0zXUFD/Dhjlr2xOG8sCEKBZ8KVNdlMhmQp
F+/33cldkWLL9alqlHGUIhfaVm93Fhp+xvmoEvDeUDtwHWqTS8OUGlsgGXRJixxO
gNqOPNiEmeq20wa8KSwvywrEN5chUJjwEqhqNe65lRW6/TwkwaaH0Jm/0D50eV9h
YJLGtEgFm6XOSmb4kJqqpN2eczmRAXus/kPi0oqEGflc/EcU7QNrwe6WV5EsQJkX
feIqjSiLwd3eNpjPoJxuuRWflDI1Efy6+NwKtaIdRBNU2wtFhZczlMN83cIDulAS
L7xUo999IVe2yQw2Es6lCvvVy7byBFbnvIWwgGlYQl8qQLWP5lNCxKgTeSe06mNH
rMGDwqg8kfgckajLo0nx3HIM0A+SoId7oxUbEjVeHhAuVYiOms2Oc4otfYKGlOVd
aE9iOW0WauYU3TZaZXDRp6Pm893DhLxpRexMpoWXlt9WyhlXEcXvA2DuAa8vPelQ
ItlwIn5sAB4Jd9hTq7vPsESOF50jIocuwx6DsjMGxV7fQUwFsZbL6DVrO7o5ux/B
gxxJZ9g2Q/PkjR9jh5DktSB5Vxr0af/c7N6lKyzPAFN0240xWAB10+MzvPyTHoZ+
Cgm2wFGB22dwrZg5aKaLp3vnUD9rpP0yn6nFS6ntM7/QdSOXRhlkywzW9BVLJPgG
MZCPiLoG5/KRXgJ9CzmRyh6Z2+aFlZQhCWhXscIHXhTFqhE66TtXWT0i54QV6y+8
og+Z7sfGb/xf+zJYoEArRG8oVfiPNyL3sx73atBfMOCmprqKmD0MWTnsj5ldIZuZ
GfJtvI/WSRgAh4PpcNxbb6bNfpFUPdkWZ2gIlyK8J0wLJ4of7q2dgXUKbCbUAxOq
c1h6Irlyo5ybjqU6E61AXJG9rDEw1HKNY9CGanwGaRXiPiNo7K0aKrYDfu4FEPYb
D/uSBZjzMZ2/hYkL7EExw5bhwtze1iTxFJ6jyzVl/AC+OlilkDfy7T8tJTz7Zs04
FhQ1wMkjKjHhDqQVoUGZTpmAsr5sBM+naxyrPjQzMw5+Yrj0VKBois1jLGHkctFN
SuacuMGYI0smTnQCtbFLJ8b300DxFXFy3D3iWSFEC3ZsomvwzbnPOtlIG+bw/cxo
yRRWz7MmtuWoJcEL9XUoDKKFSTYJziPhNoE0shRWzzuP8ZSm4c6QMF6Vk7OuK9l3
/QeUgrqFDQD6dklQIskaLiQ561zIuM18Ms0mFWsCzRIzC541PUzRy7FwlV8as+le
2fX0lyipmdeY/JMtMbxpCIlP13o8M8yWN78oX5mItrvQViyQvhAoj9D18hglJR34
W4uw+kF0VexcWnXEJH6cJulMph5hcS6UozXrEB8K+KhjmfNrraTyL+3vbtPpKj2G
2qPDNVVxSXH7wWelm0vuXqR0M2r/6Y13ruYiX1k6OKC6a0TtgOsLRnDyG9KaL2jX
O9yJ96uSDjQzFwRjXo8XbKOSxyAngUyoTFkeaO+DMMwEb6wxEv3WvmKAINgk+wBB
wy4tUWkNSKGq2r84hFyPCT+62DZdeVgGQB8i3sISKcdEJpMQ8lxA75nt7Vr2xVWt
re7s+vJru7OxetYQJ3PlceZ0zEOCvf8y4oTMUzWBvoImAVSPAP5QHJdpW2T2x0wj
TGBzSAPFHfDUhWaGBnmwQeVUkG7YEiBtc5IU2DuDmklbjdJfmIDp0ovamjiVyE5+
Iar4lPh6wrNVSbBMYB3NDg1W65isJVzEFsGWZZLylksbXoi2vEPJcRKjt5Inhlvs
OvvcFtBXfrblaNZEGV1+UvIOmQRxKfQfnyu9O9KbefDL8/p16YBKdogVO1Ovmz8+
IaBWahHfqlTLg0RJpXzofscPRT3wGjhM1Lq4gTO7GMDKXyLL+g3Cg8pp1wspxpcB
cFwpYdgAys2LjS5o2B5CR8p/E9yeWZ/BLX42ZyhToFJGXWvTv9X1Wf5AODiQrUen
3daMLZn50UQcVbv3e3ysQ0hPK6yiXFm4L/pcmeH/cFboc13G88Y9Vx/T8rl9kEDR
Z3yiCT26T5TrxwB4P1DfgiiuIczdezlWW7Yzr4KGaV/OAbK9B3yLYQ6Wi8Ro9A4S
SPxrd02dHa56XiyWpJr2eT3TQd3I8NGlN5qpABYbm8L2oZeeulpesgIv2ixTfzTf
48vsGPCmHY0gq/RJX7lNU7bF1RPDAU0coLm3T/yYkNashWxpUeIY2tSSb9aTrB/f
WUM7suZxXmyrXiEkjNgjjpEV8qMn+Ps/GXfQrwgVer7/5BBIfCN2vbG47/vWVKBB
78qixkzhowaAIqoEmPZ0P5ZThLSJDaJZikK8msKfixl2P3LPdk8QfJz135LO195M
ufyXS0UU5he8XiBF2kIlteHiDHPpomT+ypE2POgnVJiOl4XsYGQFiCywjfe3KTRg
0jQmlQ1XGSS/QrEVxiYa4GPPbSxQ/ItDvuHi3TeFah2wdT+sON2hPgd7E/zRADKe
sGaPzkpWbiabqUy6zqNp9JOjKzBV4VMkKwHP4D6/5AJbcsLj7Gdzv1BvJLEpMGsd
FrXMaCnrKI/NswRNvmabqcNTl2+wL1q2K5d8NRUra/s2znSUC30jqyeOMAmVQqoF
VVUg5t/G8PnA0BMhjqBdwiN1UXDmZGrgtbp7p04WXX6bVntSPhAwEQW4gSQ/+3jj
7hhKW6LEp3zn4eV/SurZHrowRn1CDykxT7S01ucfrqtBY4t6UBQ0K25H8Fa77V7Z
ghDlIwT4i0f65+eVJX3bxvscE4F/7zZs/gl/83NrDuNVr99L9jBhUWIYbBbcvkOc
MkqDYEyQM7Ig3hIuepM9rXLApAiZH67NMqtAt5BsR/HsMW+poWwYADvnzRrc8yCg
FxJCnArY/iYsHXWE+uhPUE9Dd/e+qcLZd6HSvZ98vY94rHKqwKKjr6qnV+A/pQ8a
d+a2JchiSK+8b/lLOs7NFedQ+aG1dXk6RqsIFT3kVEB1o0p1E6KrueKsDBz3p29g
Fyw7X84Ixjn01OunpbTHO+dokRjuInULuaJEsF9uYijaWxTKC/gY5kwZsdp04sIm
5mP8RutChEgPD3tH04nXHP5ZDTh/XImT691XjD3vqdNlG873TOvGojjxrSCe5aNl
5fkp8fDoGTacq/nkAywvVKG6qVEwf4VPsEJcQkNJ70mCK842MwT7IQJ0bGwarCHE
k1X+Ex8IX/EkhgN0UtD9dZo7QZbKNxRIJNy7OqVy+t51u/8z8J86gbwYIcnqWn0t
PJspjPRUTMWEx7DuSWXIFyTf5rfb2Kl4m9fMyYFZeVquWGojy1domD5arYWR2INi
6jz1jx6PCf2jEi5gQPE1mzg+95Yk7lWScFTLYD6ZVmMc+j48J9ZmJt7K3t1mM/uL
nKf+7STR+1OFG+UvOIxWYzTtjjrVBR4Z37hu1om8cLJddv8VQ7OvPwq4gcFJlt6q
Pu+/c1ncUeG35iVe67SaG1D1ZBxjTY5CkqUCOfNrfZZ20v0C3kpNDb0cOlW/c8lI
Dg/R78aGOgGXCwv8amYBXXC4kvmIOrOMgB191X6vGvAvNae+haRzQ6tCG1/48wwT
TtKQgZw/DEQY6XJsUoxoxpdqH6YfwJbFPGPyfeWIhlI9i4wgwrLhcVBL6rnBiu42
frbRoyEZn04y2nOCmzV6Pk5qMgqFB0NpS2iBN39zQTxZA5EzU2a7jpjUk+bj6ajf
jnm/JAorlTgdN9wDWyIVQxcnaVOh/lLsVJmlAP4eg14JG/cAq23TewvGI2NEpCCz
hzFuqeYhRkhd4JfFFW9uxmUVzhAhQRjHSmw5gxKpL7zMlWOuLL3CJmumAOx7T+gC
MDKmmI/aSsPPZQ6plcOf7fzFl0rVGno8G01Tr76J2M55NaDVUpLfRLslyGv+/nEF
P6VGpiEiusRaYj63hNuMVP6kiz53r50DJacWLOXFlTsomyrZgzFdTdklCWR96eWr
vKaUl69pnkLqFnTZlX1szTpSlzLncqAxdMB5qjQ76MRdihgqJU0kfsJOLMl5mhER
x8HqPgf5zwJ5jxc2E2U5xHkeUndfQHPLMpPMja6Fbzr01ax3EvXqbSiMbn8cu6u8
F78qw9EhyuBg4OHH9vvBBqAjH5C5KK2ONYcIjE8zT+81Vtcs+7lm6IA7zXNSSDwC
8cHOgObb5NUfhYp2QldDIUALTPOVfEQ37fNy0jaa7dRe7eYlqwzL5EQdtzd2QvDm
kPlIcgZ1ays98zvgexV+b/Cz1mawVfH+2UH0/xUjOhRCJLBEKsp37xnVENtUd7GL
IfIEQEp4quKQS8TT+pqFsQYmgp7woWJSSB5FcqA2ac7oh01fhnOdHzShQg3t/8fx
978kdu4XggRN+odNa1BtxhFZ34h6cyJwaQdv7ZOLE+cR883UFlioq1Urct1fUrv4
c8Vgq2jOo1pH8EN/I7j9YP5jDMviqyhLVUw4CDQnuVHDmfGf2fgzHR5zgwrinxxd
UTgUdBNnM/vzQctryuZTXiyzyGMTUMnm10CVXUE588/KUm7OIg/sPlXpoOz/B+Zn
4oB3pLIHvFENcpfgZS5taWdXujr+H2/Wca5o9GdE4zJ7iW+ga6cGjJmjEItJZ8JC
YOFCXp/mnMIr6g+wvKZyhLnlsfdyLggjUaXpmGoXB4P9MJ2Y6DTDJFuEMyIGaaM7
dlqQmx6nvH1seO+k9SBYheLiXbJkZSk4T7AlebPzVhnBFhnetsaZa4SbA5CjhMwg
9F8m43t0sO4ATO2Q/NI62Mg/qtCuLBMqg7d5WDwx5sPa9LsqsM2Effbl8doAQE3E
toDoTFyNDPF9DafMWB9TwKVu2m5T2S3EcCsNn1svvD3mWYcqPU8IzfxRQJ+uSDZB
IQMwxDc05rIgNbaT9L/RBwDmDujenGOOUMur+a3DZn0A9H69OSn7h8LrISty6EDQ
c9dXEJz0/uHikQ/3tGXQ2sU7skptSAQoCAjdmu4tLaJ7hUWZXiUvjER4n+aicLHm
7mJ4a9GrM/MgUQRgjcc/C1NVroKN2rK1SskSh2IZBsMN4P6JlvJQjy3t3IjzJ7hz
nl8XEzNuWxfW+wspizdnO6y2B2jEypo7KHGNM0CQoJ9TuoF2f3+G3OtGo88h+leQ
K/Qzc58Otr+ZJI4vp1qqzlGIObkuNuV0HYDLyU2P50YGbBHuYBqrEp1Qvx25x6+9
L+UNClA/eFKuTprcLs1LwMKvhAMDQZW6orFNC+LMthv5PLRYSBpD+yk7ZdtuqlpJ
TV9Q2h9h53dFMYwMv1jPOBXUA9kxWxAXQp/nZXuHpTRnbOyKOeifYnYKnz948Pwm
LNjiq8tF6VBRfxO5+blm7wom7ZEFq+SXpPppPfoXpIihm/bwCx52hREEN07VNHVB
B3Ln9VVgiqR5IyUTMnZUBWggLgEQz1Xqeg+ThMJKn32iRl1d9vfnJzXweI1Ceuty
vJtid7RNPx5Cq2PBnajiPfeBh3kAzDVN1MisHncxz57O0VUQEMJwtrPlFg8wLi0Z
BvmSLo7yXHY/V3QMmMkoaltENvcK4RiwxegRNt3r2DCije09+poSwDc5879/BjjL
7MUIGetsnmP5sUQhzUemG2PKtSkuT3Flz/A9JPVy4eShw0oBkSJPNBwizdB32uTh
XmneuVuXlGyDgRtkSjmtsftsbkEq5TXhn7hg2vFeytmOu/+e5bfmjwOHQFFY34sw
vKHqQ1N7+68nH9YfbmsrIN4PcNWHsSwJumQPODVtdRj5LR4fQ2HNXNtwL6IR5Jyn
7m4sCmpqFFILyB3gtWJWubs7+byFC9VZqg2jjMiS1ES/BWsW1dnKRdrvw6FxVS4N
QuIkUBsHAXNDlAO9e8x0It1dXxqx8NFhAQU+YiF3tgruZu7BckEhtaJUn2R6kCik
A65L6pOeSpEtNAQZjNhQVuuA4OnG4V0HsJWukDVhdKvTsH4TKuCNpHC5i+BlNbA4
mzqOTdyFrRSdPXie2M0n7QiBOrZN8Rz8j6YZp9upKLaqnJmnM6hoibh0j3ONN8mh
mdB7YX6kltq6v+Cua2ZMJOL0jeBTflBonOE7zmxF6fz67+OZIyuR1DJwua71BAq4
a/2iQNyQD+AwbqPVx3JnklUPe/e4gB5IY+sK8bRTNQANr3zkp82+sfJDRejXhIvY
4awYTEDEQDsq2XmI4FL5APTN2uQWTx/LuAjqvPlum9h/PGkWyIVgX3A3KuOlWOF8
j4J1QIbGta79IOXgeW9rDfoHcAQITG8kRtmyV0adtgYOrM7moct1ocip2wMOyWWx
34p59lRYnEY/X+ZMNQ+A7lnhOq6ijZKg0HcLGLGV41lqNjz5ihndyQ3H8RnHPGUN
JrXlwzdEtza28Jx4b7oBaMeh+HVZ7rctI0z547oGcsTZIj7dClypWpTFdR7Zwl/4
yXz+k6tNJD+BvMQmjBwSNDnOkTGVZxs/zKrk957H/nEcd/z+ptuWym9NZ+5tH+Y5
vZmnRYVplXCHgVkqrMlNoh4dRXegJvqMmoOiN3+VFZtKEBiOrNKF14mxadEfTZj1
p3NVXZMH4BsoUq9ra8g7YvGFC9x2zUpAOeOkHyGJ02cdmyGKR0cMCSP2kZJgtvug
kKWxJCCqAxhrbZEFgZIGYAuJmTSHPg+0HtdmrOvnPNKJkejdvYMB0sLG54HJJ8uG
VFCsm6YTQ1B/K6SFko802BlCyvRj0X/VOmuZrpvAP/fpXdzL0EpVxsCnE+u58Eb+
KzffAy8/NqmdpJZ30m9B9HsEqV3FakA0U344bESSFD02mtuqOvhyKTE5yyLq52HP
MkwBZ8v7Po3bl4P6ovKt3a0LeOlnXeTEWX69sURGY2J+c5+YMGWanuLDcsjZkH7i
Nc39CPxzu1zJ55w/OsYX0ln2Qqv7AFcwYNU/hdx6RqZiUojvShTmpo2AtmC2/BnG
rdf6lOELDSmGpmRlkFbvKuvTqIMl8N9/LsZTUfQBeLQ/UnyLeb6YJcBCVLuqjryF
Z07MqQeexFOGn9ew/3w6lHblW7Z6Xo+5+li6D290ElP+reP/aJOygE+MGFdFySKH
+VAzu/OFJnRPJGbeBVwPKfL2C++qCHkTgtKqsNCQFU7BxwQJmE975a3tECGTiKbA
o+zFx1nAHiyIdbi5GvUreShfsEZVGfcFVraxRd0Z3kpF0+VniUuoHslM5gHcRuqd
H68uG8D8cCzs4qnhHSUzDinghaSPj/tPadddCKosFdMW2k/lOcKLZ33+oq4ptUcv
L/47slE//Hc214JmsVOmiE1F718R05+ZvSI+AfpPqC5HA+hnK4mULEkMpgcm6UqB
1JB1VsAJ7rqfOcgHuVHUfghuPCcQ3ugpFg3D+tQuxciTWKvs4pZ0FiCfzb9D75T7
FEpF9qJvrNlCyeNBoiKauVLuKcQ2c0nOvyChToXPqkraxLVJboF8Qd/5mvfl6G2q
8gwrmn2jZkxaExyaOaavbvg7txZUvqo5or3aXkC6Cv2n/SzzWp3DZnfwJy5wRIBa
2PswWoS3tmV0l1XLsII74vXSDqwpts8ynVVjkVp+UiEFlrEoM0tMQRohsiiLInF6
D8MeTxyVDbNFbuLp7bl6pQLMj9k5NqDawzUFchMnv46d0IeBtZ3A0acozXexytzS
07CqKXIo5Bn7vKM151JqtT2/TvfXgjrra9Psi76Kd3Ds1BiSX+UBLBcubofNeVSA
+cE0DtgbT8Rxfwpq6CYpTvrNmzW1O2OfYKJ1/KmvcOjCXPdfUxxo7gxN8wsK1zEN
YG5nwB4wh27xi54xwP5hCpGBjS3clRd+IUgvkltzfs1IG4ggw1z0ZX1l7rT3TIJq
xB3es8tNkNr3eQ50Y4QvMPIoWkSCVXC54/CbNthO5C1mtLnIJiRgvcbK3lxI/caY
ewtOSEzpjX82U2WMUeAxdHe/Yplg7BzcsMkcVKsOh9/cvUP/5BwhQC0UABz49R5n
fGKAGHR0buGAhE3N0oxV4m1a7zgxw0BWl+uBxdZgRFblt4PI3fqdHuK8Xp0cxNL2
EkoqOn+p0qgdvAO9R5aJ+Qv8ai9FZjdEwmgqutd+leoODoPH1lQQsKMdU15SP+Vs
g3fdax2joogNXK/HuA33hG9r7oaeIWTaINWfU0ZrO17+JhNDncNzsKXEwxHxHoPB
DSh0q+LXYe2aPmJXqvkRpoNKiQsDusR+czY23hJl/Gwb8YI/x4zbfMSsSU+8mk3G
Spds7onrcZA1u1vDdNOT+0lWiWSI4M5GlWALjtB5MgkdD2EQVYUrIuax9uMFi1bl
5EnofRuYP3du78UvCK9pLk9dzeRUh+bm+HrJOTFIw0uUAwwp4eBaIBO6CuK56+ed
G6aoW6ES/a0CizKYHQOx7qd+vST75efuu7h84h7sFxtAakTapmTqaizwNO473laV
uJ12+z660/mQWp1q1zUeus5KOuq6iQbwZq6aF6TwIu57T2FMyPxPamcZw+b6nrJj
DPJL6OL8ll6q6XFKfzH1B/Up7NeZj98EVAYPZsJi5BkdY0hlsQNM/VKWh5/PneDe
04DVPq31DMumOSHMYo7HbzOjNXiZpFIyOr1kcPPIjPBwm3BADJyi39xATJncfXaG
ChtoGaVOyXeUP+QpZGbGJlQpq7fcB2rz+Vb/yXw3OAMeFR266p9AnAUtF0E6r7Qz
FLMJouoRF5MAj6CoHiDO2z3RJiTNr+gQd6Qz0tshaY4iLDtHNREBWec72853mDf1
ayu1NHw80mYXiO28Bqos/L2bhta4lmQjbwSsGvTm/AvP6aqLxlvIJ/jQtIxWjZvk
dZZjbbHCL1Bd9IXIE11oHZa6OeGW0XWYKVYaesRx/eoTn51QfN2QtJScVXwV20Iq
HC1zyrgpOesCXDybShWs8fIXT1stoNks1hykRzuDkBJvREe0TARl3eZb4yhJXZha
ay+1ubHhURp/HZdOQ/Zf//4b+ETSoFyW80sTDQETL9YR91YyVaXAIDs0TSHW2Nyl
694+IFJdR1h/EPeS+tcZL5G+wKaYTJne1yRvsSrzv0L4HHqgB40iZm3HguZruVYJ
dhQjlFqLqASmAcvrZsUzegV1LsgiTr4bBSV7El+JRLLUDx48gPgRCIn+A4vyQfo2
bbRjZblx9dnfIDHLXpX4VBtvhfrLsD08rQAIsmNBx3XvSD8pHkvPn79qzLUeQZdW
ZThO1cTvOBFb2gxb0lYyV0zS8ExFvVLOUNe8gZte9osp4pESA0KIrGZJZgI8K7Ju
LZIsc7Ix2T/B+ckkqOrGllKbO4m3EN4flYRZlVPcuBsKgEJ0HefYJ3Mk8r6HLqtv
dOtmok2OCzNh2MzqIGbJDKsYovZFVCXL8t4VTWaeeO5sDLU2ddVCWyTYi9pPA+M0
HdWaXd4qfaHRnKi2Z8kYNOcptyVtI2og+Ly/E0K+ybTSRo0p+OF+akgGs0jFQp4b
IwWT6uDAFJwEkjCp/JltRp8oDvBUJNtr995p+t4aJ87kStYPqhjBbo84BAHk3bRe
7H2kx5AJ686BEeVexK0CzxP9aXGiNdalXIHNRd18j8O3RocPWTIowmIJVwKgYCAC
C3njZp66e4u9Q/CKwzPn8EfzWznDx+uuj/CH5JBW0SPRAFZYX4kdeblfOlHMsYB8
znBCPubJ7XHDcTiSL08BExWYFa9GvnfBRRwTYk9SFFO1Oh3X+0hDj9Yi7fD7JHwZ
HjTZ7ahGNiDB8ri8WI0x61QvpoLi4KZY600S+RhNVtatlGeOeCX2NqLMY4I91oFe
zLwoMYLUrqDkbRotBNgsUgqul580SEkBPmljBnNMx9Ijcg9mcBbgJL4CjYsuL6zm
2pDvCpNywgRCnO/6QYxpVRGwWxmTwF1qldL3u8r4sSEIjOSeWTF87/4CUg6Spvcy
Buftu95Z6kjNSjbOwJAPK/aScs2MmPiBCCtiOk4y8Zt9qevExEXkJC497EGCDjqh
ZA7ZERQeH/igCaNf+w8xnWFCDtwBIYqS+bVz1mN/fIrPiNI2y8IzJY6XaHeIr1E5
17YTJ74qfCACaPBr7VLYXxtZoWeTlfdHnxbJ9nX64ba5HTS262ZN7lh4CYRh3Gft
5fPMsnoxstHmh9OW27rhoE3WRJKVZbjeAfZqdmK03KMf1sUNzwra8rR1bcC0SoEm
TxoA2W8ZWkP/I2uMIbuublhOqPHZR1GVPBXjVcPfpT8ktCMj2qacTgXRix98NXAN
2kNrPEAxM+2H1Mn7TPNiZW+/kix9Y3Y8Q7eDOo/uI8SZTtTjsqrfnZGA63fd37Nu
6IA+Spn1Y85bQu6BmCuEdNIQwn/ZEhhD2Th/3gLDiFabt6xZkqCS/aGtO+Hvqn++
LKPiFiMmP3aWeDukZns1PxOgyCpB/iqIZkpgzxHoab8h5812AcerMocRDqevNnaE
LZMPxqASQfVJvzkIbTHBOwazozgHtvmMwYgv++8G84jvOxVFt8riCezqxN+diuzE
Ha3fQUWFZCELkdoiXfj7GQt0Er6aQzzp+MhxjuUwU5sZxmhgl7TmqgDpdrMKR/2j
QCYPjezU3grd2+nP1mzMjT3Gfz4UsS8pXHWmsJy9r6Gqs9iwVpaoE89PIU2a2Bxi
+F6YNPlYTCXGXG72NBjCaEoptT3v2PE24+vObMEyW4tb6uR6FSCnXfutZffN4TSL
BuAN6Xav1Fnqs5y2suk7MK2o1wpzH8+Jahyc/riNCWhB9diXVQkh5W/SAwhfCmqx
kCWmgEeOmBPRvBqg9rltC97DQ7OD+62hlComfJNBDKcvh48bNYZIfxqgi4OvdIcJ
EWBy07QqtyP3IglVbUppghH2z++ouRfRR/j/MDivc4LZwOmpzkoQHa/v3eF3nB4V
SSwzQHTfeFN719NJM49I+DT6FyRReIECWpVDqZsHsvlK8CpBmk++iXZHmhHJQlJ4
aNhBs4sToHQZpgAaelUgbvZoQk+LekBcw65RairUgPacqkvuGj4pudgQQTTJKBZb
F21e2e+nJnSNt21hSgVlF/YiE41mVYJND/eHuXdHap2cFN7mnjKwA8rXmWa/jKiM
gsKRz8fNfQy12RKefOUfWNPPS3VxsYjyEwkTvcmkh/SjKco1ONKN2HobAkE85531
lkRexsZ4uTuYIzwKSEhh0OBZIqDO1KtVxkGNwQvv3IsFiBQsj/Vz/xM0zvU3DT7J
IrqRhP1c8sJWqnWlv3V4WgyYF7kwn7VcHjEI9LYC6tvgtgm+FK/9UI3J9poIZfqO
EoPBz9RV1S2zCNeXrWSGi9WqsOmP6Ba1rKJCBfyAsLV6JNroUX+YM+pOpNcvhrP7
tduiZcTmznsQObrzun2zNOAY97wADzXZAMPrgBpgkt0zCs/or/DTtYxW5iv5EIMn
I+mtaNZMi+IydciEha4fRE/sdlERP7WBxcAsCIsANUggASWTLVsjWrvJDLULtyjz
L/CTM5Turvjp6EuLW1PDdZzzibL82rllrTE+Yg2VtX6/d6Ohh0oYZx8FtbYX107V
jEp7cHKVnhcWwO2+66NOZZwXwcqig6IPri/c7eJwGwEohWJznMShj2ev5pwofvpr
X96a4HurMqVVJ53L+A3QqBO8eUrpBY+OFI6hHThSpsUwIcnDORwovspkz7FhAWPm
augsyq/xVPshs6xSRwpMLu3dcwXQdMAf1SeHeHM0XfrUfc4I32LITisUPD6TI969
bvb9W/8kqlMcva/bmh22gqO94aTjMfx+JnHSyiOt0CgWDMrxAiyKZrharwiyMq5c
2fx8FuUVWC6F5nxLZoVujWAVXNIm4OLfcxhMZsnmOmF6oZIn8t8lME8aSVygOZ+M
iBsoF8wSlq3BsgUZuAF7WT7W9iDnyp1bob4im6ffk8cRsR3IgyvO1f+tClr3kmdM
h3SRvdCLJkt/IAEY2dK+Y5aLGXhY8jZUGObvIHE5u6EK7RGl5qo/AnPOzn5vxXxR
1Uqbw4oIUWghR18/UVbTRz0a44LlFcqfilYvU/IQJ47g6yyBpAVwE7LzRK0/MxD9
O/dbCVpojewB1u3mT6/aqtb81ay5R9UNLI0mttQYePvv25Mw1AYMYRSVp8XGtsUx
CTwQJDIog7C526RpcamJh84Zmqr6FsJO6uArkjyw8AOAfUf0gRUbwG2rtGRFQdVU
OTCw+dMDOzT6fZ1ZBmaGpsE9FXA5TN6Uum8ze0EZhOGS/Sf0ZzGNbEovWKCvS5Mt
20ZO3bwrVDOkrFJxvnnA6qWw0EM8Cys+GhF4f4DSFfHytrElAxY8DHoqfTL2uGtv
fTUWCScAq3IB6GUyg4IAwIMKh1I3iXv/iF1bzDsTSpuM3ZPW1j+ejyTwHmdm3M6e
kwqtuDkBqMc3G4tDdTOMeMtzeUxj/pA4GuyF7A7UkduVuGfxxXJfJl/HkHc049gU
ShwDZyKypGFlSO0lHVBCUGlnjWWZunl4yjLTczvByXUNDF1DdtlLPI+K+Zw0oEs1
75eftL26ISiW7ZjBX3M6ADwsIpBvwxzaeJ6Su9morg26n+liNiP2m15ff6i6qYCF
NAWdeFAUeXumJUkPbQOkYTyXMt/wtnPjy/BcuRe4mgGWsuwQ3gjGJSxTuJhp+k3S
A0cRhDJ3q1590bJh4K79aB52aG0ac2Org73sIs7pAT6QsxNguwas6m8QbRpKNZbQ
lZsnzvq7KaYDmqdZv5Rjv2fxoZq3Z+L9qVC7QP4/T+x5aJQSFo3VkAYBtzsxW4dh
LPpkrNGwz01aetI/jCXUK8XXiqnQu5B0WYXf4M9dx7AZj13UTU5QDiPb2vW5uAz4
hPjcCOEtivdwtUNZlkQbqGPKZg5gC/qIAMhSWvnZzDm7BnFB+cgSdBtObxVCltK+
1XlMo+AVoJB//NTGCbK1/0Bvv05pQmAlhZM6Ap52JJYyq3GcNXUA3Gpswr5Rj/nh
yuk3SeGEccPUZd0cDzt1KYkR6UOtAwvcnhOZlMTXfGsgdOY0Gp70dWLdxP1fAO9k
H+AUAbrt3XUmOVuVFDdoJyIfGCHz2dQ/28abkSjiBUpF2GKnmur39ipnQaJ0Flzw
QI000NSbLtA/ZCi/ThPbNctPVl4Ac3Sfv2LZ3+N+614FyIHN02i3c5k1XT8FlDEV
B5Roo8TsoMFQ4+tIiEfC2Kvn5b4zMSThyftWGLduPozdAQ+B5ueyEwY9LdK4ptCL
I522VzqjECOwPWDybGDMAkRpjoq5z4JoEHBm692vuXTXkzaWlQXRzHZ89pzzLoKU
RyzgGBqyt6wwoQEoHKaK3NdbMjyeRmVtfxAQ7kR9d6brfej7Z9oJ08nV/1j7AKL7
iPmOvecShZJRvfTJHvNijHH3MfY39ckqYH+vTCFBe1AuPBdLWCCHbzJX5HgwFQSP
0qqtzAVgu3QR0LIOf0UUYC9vMVQEFlDyfxkn38DTFasg9HDLXOPF5Vxm8u7BOpov
goo8OF/CwH+luAfit28yMPAiSQA651yyfNLhi9o/fNalK7n3AiK9DAPQ0j+03hI0
17mx6JvGXKTd+wYMkgmgkSw58ngEe1uZNhOFo8NGvBrQHlrqBgsiuPry6TB1PAGG
1bvSVqFSA3VbW0Nqoi66ZRuKJ8Z8rC7/V+YCm46R0WNFxYY1Qhin3X5l7jhjlNFx
933KWg4jY9C2vSfFD4GPFwuh0jshaa4jvLibXOqT8gQ3UCi0PaOUrjGdJW1JkwCJ
Sm0hbU8S6UttRB0szKtO2lJHpPGczWVaEp28Ej/BlwOwpNXQlKzrJFMrd5t1HCTF
qRHi+EI70zUedYqUhhtC8TIuIReAmg2wKpSzMsSw9EWbrsm5dS+0UaoNC+Wl1tt2
teZa9no5sL4MhS/HYzwZ7lU9E+AbyklObkif2HbJqNIN3dZ74nVAiCUZgXB/+pQb
0knfg9EwAmkHh3c3P+EP1RuhCrzzkxkhWVcm6o3/TqMV7S+clLG4chYfaWjhHYCX
gjONO+OHM0IliYi3lnIDCmoziefnO2t58qRigys6X5G2460+CC5Zn6h1QXejaayc
1pS7wQ1huz12d5qakTuNsVy+YB3NDdu2GBvHfYNZra5ZwTvqqqZU4rExWWSZt2Zc
pAWArSRVJXU8oeuPPGvX1/E75PcVcj8BwQricmtx9TUPiVbgsoKxYHIyIZAV2uMq
58q79CSux4B9TrUTK6d8UD++f/FPrnivEmntsrYJR6xmxwWAqIbrPKQi9XOKz4LB
aE07DShdWSANnR+ks8zV1tavYNGmh8kJHTkVJq6KevockX9cmLehAFsvjp9vG2w8
ckNtskE+YrilD8QCo/3MgAltBVi7YRe4AXe7yVI6lCWyaHFOS6gm2bMw8jw0c7iN
51A5LV9KRy+tXaKXdcXSDPSBsGWvzjGSuF5J5/1NpMF0Irm1sMaZstbpOhEyu6oW
jtrMlDMTmCImVmKXo2Edo2XO79I671pqSx8REWQtRG03zrB0zNC8RuRVcLWE0sks
FF2r3F++EbRhBmmVhZ1K3N0gRlmXn3zKnDNh3oofjM/TQfjxSonMCtB6uw3DaQcf
5EjZJ+iDghrKJHQLM7DXiBXACF6e4cc50+wOvUe4iP+GBNIcEKHA0PPU6AdT8+Yi
IBFvXaBnXiNKEXQpz7zbKlnvosRnA+2dSdrn+v9OtWC44gmfJL9hhMXioa2OflXZ
dit3bIady1iHHGBuuFZynlfFzIKAz5cEG1RLUGMq5jkgIfkalzV+o3jxlmFm05u6
HfIIC7K4NaZ2UFYuwnVnOBPJpVlwK/vG+GgBA7SUoMoonQnskOr53aRxZRSed//k
wQsPw4qTCGrfBrZqi+qB73fDFW+QyC5/frQGvT1Dz2UMEJL4DqFSK77ujkoL71nK
sIW6HnaGM49ZqoqL7o1RIJ78LCtsQiUu1/IQSPav6QppqR7QAZ1+O33Kko3o/3/4
8qaxrpovja3JVYb5spbd4x1DkSAd3txqukZoZG4x40ebpVIyuAzsHTBP2bkl0qZ4
OOEkIlODZmsJ/2g+04gb48fHEUVttM4PhM3Fd7RGvLOdIH/QP2Dcbsd2QCS1qhPo
CI0SeVItAAd0T14SeUxBEwMA4fKmxZzsvjlXBCS0eYniH7fZ1iukiHy0btK0RatL
SWnj1fRO+UHYRHFo0VuJyXPwKpi8J9FcQWvV8BIXin8OKhiceN0o9atNRuor2kTV
V9fm7+tRvYFbMBNCqhHHTCFUFMUJIZKDKtjceTsmyC48W3gbzepQhC/ZnyLZr5pA
XzxkqyYtZs53MpbsWvIpEKIsGS2Eki6n+SmO3Ug2svfXjOAzr3luguL0MUapmW8i
Ephxb9RxcupBoYc5vQxPTgxgA6C/NjmIoBp9lLsL+bNfneSQqNs4LIyA6LWq2D1B
pGOj24hHnVRjJE5FHKmYUyb1JJYpTkpgwaYKyI+j6ed11uL49p5tAf/K4jXgj4Xv
6THLtml1p3OuoOv6PmhU3lXSRcA5p0ii3/KAcpXVBXhez+JfS/8kam2AQMjZy3T9
lWTjwlgB1Ma9Sle/VTGoMz4HVDU1LuwJa9h+9bai6iHFQkzI8bUU7rgkDGKmwS59
h8vTOwMFMhoIekeW389VC6LIj0XUTOEyWU7JNVrC7YjlVJ6aO12waSWpqoOdcwnV
lyiEGzPSzsrTJANOVh+9vJuBVw7KIPDZ43lyPmGjGznD8C3zrGowmfDHH3xiDrh5
tavbjKE2OIsdjs/VUOetsE6O3sOF8FTNz+NEQ7MpBYSaKcWq7K22AnK/q/xnVpeY
Ks96US73PLCHTQxIRyVCxBIP7iTxMC+UyIE0s8MiUZQkaui2kPCSPKivPps8tAsz
/9eHA/LuJ1KZ7KcOO3tOunl3nnwbTLI1Kjwc8eIcZd+kVVf308/ZG764owhKrU2M
2VbWvqm3pVFAhrkihc33KW4loUpUG+2q/4QvkzRq0ntzCfz9tbDWJGP250dJBmH/
91t0jgmp2+yukE0niy9E6JCMApLcAgEl3mH5n5HC+4xGPm6cOPgIyJ/y4Z0aS+R5
0uqZ5ZNhkupWkc2BQ2VaPhBiGXx0hPKnKgCJPeaHWuRvulhUC0AYmBBaRRhIgz8p
tIMijjqSnTA6CPO2FkldXThq8UZ5rQBmDJDn5kJ3lVHdY69t4x65lrrg7b2cPeNX
6oT6GMSea/nG4P9EsxUvVgiftC134MbsbM3Kl3P+JdofVvuH9jS2q9RmDp7ct62/
37NmQWFZ+NMgOuFBt210G/GhSsxDf1v1ivTJMXDnk/boUaWdVgYujGNEu1t2QI5J
WuIStXpg7/fCE9fmfCdGStDiPNSD7F/o3IDR2ORI0yFiMSABlqucn2Bhhx0XHRuy
kdMJw9qE89gUypDywXWPEvaWBRYI0uUU1BkpfqO1fwBW7jWvfxDY/n6bfZn1Rt97
mKsOX222bkF0tTkSvuqrf2v5k2n1nsxIsFzKOZrWaLFdoiOHthIRSCbxO7s6Psg8
VEkd+8yAOdIG648IEfVJ9s9W5989+U8Cek5oIQT9NdgxTFddFyRWndu6a+mOG30F
yL8yXOsDLcDpXOl5sCgE9fJD9Ejyl84HxPcga6rHCohLNRuoNQL113VxRT/h5P4z
FF95i1nQRwCUazEqW2Ct6V/9lb6ZqOw5c9MTqIpfzddynWPnxLEJBeQIQd2qzvnG
EiiEcF1wAyHXRodM30vQ8qPui3906uO1+kwUTwfMUFIaIqou8FCn7ZlR3WXPe6IF
00nAKJh8lA6kZW7XWgYa0KplckO9yLNT8jhk+VUD5kqt8kQ0yDYY0128kADh3I1b
5dde3oLLTDHPH9rcixAcu/S9sun7UaQXgmWRF4ETC5yrTEXYNefUFX+43N72wXny
CNsYnrkOpJtFystEOeltLeuIRygFyetGlusiI4siNPCvUgWyziLV6zO+k3no3rQ/
XFwwAutCdzIoz3+2aZPxIZmj4Q+bb2Wq7ujw08YOqJFOYWPWDVH6KOAR49+8ufcm
J7dQri2T/7uR2bP5JE9Zf8Yq4h/AG/aYVenlz79fpOJqHqEkU/DEBzG1QknxYpnE
9oRjOOljPKEXTjiVNjH++BLEp1ju4KvS1oJf42g7Wbi1cnGHs2esFE48L1zth75X
1PFCKB7RHWjaTLr0Ji2SAFkfeeKDOAJZ8r406VSkZWTwsMTPMHZqZnOYiXkI2KwT
BskNfrVqUY7J4qwOoOXU7p1oz2FloLtg8h0XRVXlAepQlU8IBlze2jJC2ztCgy0L
a/A5ZBX4LM4DJPnQErIQKYxguxouHqt7QHnQjV62o3j4RSvtkgDtHSKMPXedDftO
SN36dlYdj7RWIFJOw6Cy7sXK4/3ldZsVtWTvI1RPUrZCNvW5Qd8XG/L/1UV292JS
YZrc84LydD0WHcRT5208227dkdS7cXmdj3tWu8Ff+xVE92xpJldfkO00eDatxj19
xRgePvZCVIw8dmOFiTIBcRnQIzA0uOBp8KcNnGp7kEAf98O+fS7udV8A9PqnarGy
IhsG+RXKw50i71jYTGVfuv1mi8zPjqVnNwGvRQRRuSaDO3cUwZkCMuiy9PcLWOak
9B4+bmIIjbcr0EQoIV7TiGczhlrruiPoI05+qeMxvjPDqBOR/6EC3t7aWXTUbK9E
RZC3ttu/dwaXfMGjS9XWqOE7aBCncb9eAMQLXEiDQm/lXqFXK4Oi7PY7YlsxbgDp
pWNnzVrHT9VSeURcNyQSqoLUDblUb/xPOy8tuN6B6XyYf1NozF/iRT+BhU2/gJa3
oT3wzjp4jN6kC0136hPK4Jebx+eP4Jub6rZ3f1u0eAbkoKMGdHYBCN5fAk5/1FNs
aq2GJGJiXv1Xl+41+F2rXV+Mw7ms6squKKMQCY9o/1dhVorP7WpucZbkNDR+nGdm
Id6VOoswikh1uiloka0uvjYf+cP9BeZpSilJ5COMgDJwdXbid32fXJRARhyjCOSC
xGoZj/Cer/TGkHJaGVtsWgGFO73rZmOIEHXyzOmNUjeWBwctCtUe05Ub1INc+RRd
N8onKq5vu+DIk3Kk/b6EHdTQ06zFAalHrLvBeHQ21ll2NqBJJdm2faEeIO7R9Azp
OyYbSRfvOqa/n736G3Zq1a+CIZfG/Kawolx3kTUgU5gAiFiAM+So9l0ubhFXGoWb
hmoN3cvXqi45aGOMEnvW3tYCEdnvx8YKjRNnziz9sCkk+a59PfHyVQ43d5jVCUf0
Il+6+flOt0k4AOpEVBHoiJkMFp4RU/Oguzr2BgII7gZjlWDXoM4Kv2h4z3cqX8Rv
NUhzHyq1QuuygubJCk10NoT+I+0HbGllykyZcvZSFK4xW579GTBDp87j2JYfSeg6
5Hw+qzJc7y/59uGBQqq6UY8BmfrUzSualv7RBqlzILddnb+yL7y1SnOkLPC92bPv
zKjBjetybs1rVcyBvQYztDabhfpU4AkS1Xzy0RSXz5uVhFaZNAXHR8erVoPO/Aqe
/S6MMUMsBQ8SIlWhE7684Ssw4YpfWbVkTgsHKywx233ugbYVK73sI2eDuILLdsjM
MnAX6FhELkpTuoL3zWhsD5gBwwqvBlMnjGLWLzXGXiSnFeEI0Q5m/8fmYzW8x2me
qww8s9lPFasmDkvt5bX92BmdJL6dc6cehE3o08aNJKoNt1DIaGOWzSZc4HiFeRjl
i/F1AqZmbJSz23LRUXCb10ZMmp04N4aWNH9eNrkWdo/XYZs4UdL4Up9H1W5BH+2l
HgIWK8ZugykudROJLJQ4Ssnf/YjLjG/ZYd2CBktvVR7mtrvxCRzwlLTBw/OKlbV5
Ps0LhktI8Z6vajZCPwV9/4RBdwCjCUCpVra/rrzVaZsMC3emdU4f/A04zterxMj9
pmsyUPhDfMRIsySaf8by2Z9OhbG+8cIoPYrZO/GYcMtAst77JQn4r4Ru7rtVJVAe
q5JuQtWNC/mYjGj1mvGMdabQtoWo++aq1OAY88vJPB4yFtxG1HiebwA4M6pjBjM0
rKklzUN3PBw+Wy8gC0Ur390RzVeLmqHUQvdu6+YXSgGLliM635gSAXZJd3txbNts
PB+OescSnCCTGkNLqZPgDcqEOwYOhN07USd+Tx2waPk5j4xuRCteyM+QRE88rDtB
sWFGbWHhut7CnR4ttTRdlJjkmsiJhMvu43BT+eKkPRo+0Wbcsne3EqW8/s2h/VeQ
CXeMkY/cLDQrtvvejDSN/+M3TcQLHIEEKOQEBT/8Ug9bDgMTVCUoUWbSlIFH75pq
zZ7LbVTlAF3PVWuZF7qAb2aR/pLBKUzpAW2OGzCjG0WfTOPf7W712vqaPIMnhIad
+NLtLxzsWsJRnLcU/eaI6QA/hBhqBUahbg6HzSi9N7KJtEEa2gPHJIZDPVzyc0Oq
PE54Ie3wpGg/Yz1HnPB2jqkB86bzLIlxTuUlRGIR4wlnM6AMHy5NbLXmnQ8+joq2
7fXuFcF8QcMspCEZxH4u4WvgPo5Nqc3YidybP5Dzw9P1WgWYMq2ueRpLqATnYye+
T3T7rzFuDxr+aXSFhVzZB32mG7HZVOARhmHKohI+zGyk+x4JTM6T7oQaAbzAo9qC
afP2Mwe0Eh9wbBSdGqdnLWZ5VT1yRrWjqn5eNoL0OgeSYH3KUfuglIH2haCb8gNI
Y9ytbOtJ00oNJv3+vgvEC9JVMPTEswwNSAHqaZUEHyE6A7EaOLEC1OE2Do6YuDtK
RLFwRBH2mLsz95bHiavCCBTnEq5IzepdTw2aCQdMsLH6iVeIHR9YMYEIFp3rYLwu
sxbNBG4gSGRiBf42vhNIydYHpr1v/JBibVk8ViFk/5SH1wXI1mwRc0ObnfsEF86g
o3fiHsp3GuGA6uKheA7iSEK+EgNX06LWp5hCJ+f/6C9j6Jn3Hvp18oFCGjrQER9b
7UlTdSzlHj2XPm3iJ/nHiKXdN7xBZ2qdLmQk6q0DGbkTov0XiMldrQUC3k4/sFYw
fmLVnDHtOWmmUzNyBpFcvAqhuDtXxmNCTP5FKRfqSY5Sh9Ix/vhsu6nNWk3tzvzS
DJHNedYIbvb2aHzy0h3v6h96rIUGbtmv208HDU/+Aegg839bNHkjxMOoP2lM98O2
CrMf/0yDYd+QeC68uO/S5cdOe9jHiyaDNaqAvDSR1awQLlxwPILh1dNwJ1thYOSI
/ifG6U18R5E8JSQnVtBuXUN4uLKjnDA3f9YC3Gb2j75/gd3HYEJC7Ss/GxCmk58d
5GDHHUOd1oQDNlkhp9aBNf7og7UD5qp/xyUVgJEdtMsRfld5Cc/iqt+StF9wOfMI
eYB/+uM8jocWw74uHaDkeoQOMAdv2PiZcYnNVF59sEKGKcjyInR/JbXVxaMq9QJe
1SN+ANb7KbvEji+aQTn8ly+FP168TOuX0bThdwpdr86TkOREvX3Xd82tOM6Rt6np
anDs9d5vgdI+yfWAAlESZpltdq/YU2V/pzkr3w4+O7KvKLt3TBEtn2jO65s/uNmF
8ozLClgW+p0+9RCdfcwEXl0xajj/fA4MEaqN8dUQYnq9nyLeIZB9oS+lE2ZKlBVp
fq+p5wh9gpowx0wklcQQfYb7HeyBs/GB+pKVkAewN0gA5U8p+w17aWi2XXIBeScK
QksJTwwxuD/SVo2mcKTQtHpeo6gu1LwAqQOgCtePmIjaVJ8pKAh1+AaQasPgE5hH
vn4STGJplqb9QqASCDYAP/3poGNGScW0tC2Ctq91nEgv5rAgzcue3n514rznxEFz
bCOQzWrLM3/UyjLZS3TiH/T9t/2/KaGecaAQ+9UcvIXYr5cSfqW3q5xDrtMqfq0f
kY/XpA1CTAHshKkhwymwr0x9PFDocBPSGJE/W68L187Dhi4A7mxiVb4LIaibglRM
ek+7jAT+ER2wMwN7QQiM3LeLyEScojP67UzzGQK7oetYfjhaJ8eOZfFCtn+Jis1A
YsG/iEFXPohNFTNdkgiuQV/mRh9FkM4fxBmgNQ8R+lYg5zuzaMHmk63RQN6BHs1C
uHlQtYLK4UmHtFNqUn3+Ih5lcv50KOV4iR3iuUzd7ITK1VUvBGRP42azX791ZRR+
sx8D4uLRwkwvfmNUdjZIvU+ZhXlgZxEH4qnSyTlPxzMfuZ82wDEUbpQIsZ1gbMy1
1G/F8poUHmLy7b07yEQxbWwG51Lmy2hBT4QR2ySw7OE5Rpm/pJrS4kEC+fPVEH/D
ib1PT7wkabrhzUBdVNPq5XadXZX2VUZ7B1XXWYy8cVNvL52/kjWoh6HwbOmcV7kp
A6POuQyta2IISJ7EJqfNzXTd4BIzI8oz3U111marU+x2RRLwbRbmaR+DahU6ifoG
LoX/bc+YHXfMidXJoUGCfhcS/LZ8egQ4VSnnxTOnMnd+TPkC/RtPpLn+3ZOFQ1HB
FqP0JTfUUzNKlkCUJFzV1EWlK7GWkCvjAtXQ44cLHMXp0T6BIcTLcd1vTpUPk5E2
yb1tvpNBt9u0Nq2og+KPkXg9v+XO1mPrtL61GNcT2i5X6pwHYsr3Gp5euDvbe//T
KR5dxVoBJF+609Ve7zGHBu1vdQaJeFVEc2mf9Reac8rRUZ1CBlg4Mjz7gbOBLqnf
T5iJDS/e9nzCDZKW0yb7HRXqQ7g5FDu44z53yiDICvNb8ZvuMBcZFiIJKUpNBZ7+
yY6z8cJGmtBj2ypN0Bwbra1LeiYUCBnPvsSXnvp2cP16d1zFzbBp4SKieQvTotLj
AEKdn0Ogr6qLzpKzwL/fLs+wZkoa+8cpMHkwQeHEWunTcFo/z7bIgZ1f93JzlYG2
WaJuQ7YefIdYZIlwX76kFeiP5ueGtlaUoKUqOufSFpUYAaSHcF0ST7WG8OS8iX5m
`protect end_protected