`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1648 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
YachDS4bpHRDzLXFQC4CtUC/J5nUtBL8dlqNOiLWMaKUkurgirQ+/gh+DEvpf2K9
UEyI6SOOfwqcQy5I71DyU0QkvIZvuUVdBxEiWm4pC3OfRjTN3swo4sbUQSPYa28t
Dv0yKFQ73DgLg26dwGkCN8CJjTkkbcYiMCUR4mvakH7LkeEm5d0i89g943QYxvtz
x/uJwZfVQd9/+M+kHxdNBeAEvNOsadPwxehFHkv4zD6U8nBaoW1HN5vI9Mm39Kwp
ZVBiEa/N/t58i6CcC2U1hsxTWzBbqJ/BX++OiqYS8864kezafNOE9zF2zw16uMFc
irzTOr60wXKbxDPTpbcSuOM3XVpm1isXRv2P44vAsvHSyYZAsMvzZFCv8m9/1S7M
2ed+1LXlwxyFyv7wT/QS9t8agWSqin28MmWZmdsxK/5/gyjO0P7MSILUVeP5PR9d
ZLM0xGRHccajN/xtmCrjG+0uuqUdXDT3W/oV1R8xNQncKdBuLYKRLAW3Hfuezx/i
cNW/5PyIwPMqeRGDIlqi1/qpRTMZ4DvpJjjg9QgCkZ1zC1AsChhorJWTLRaxix1Q
yN18k625nOI1UWGVVwO5I+Fq9jJGeb+7CcAJgyv4YzjvsCWMJj5h8CM1KcLxkMnQ
bivkBfrzEFaOdqydCMe2OB98gNeLYIyZVtpSplOxH6sYxAYCCI1CCNHhVCONhYdl
BdEuPwoVuK1nLGCQ3B/txJPAQzGvM+rzI10VYLeDHueX0RMj6B0YxHtCSfdd+smk
5gnwEJx8pZQEHRwj1W1cqWlnnJ0YMOqvjDmXeXDsavD6/ib4pLKDzeOC8THCu3zj
2ABoaN07SzQnXkkDGe28FIdg3lRKW+bnxr5wWaUkKcxlgUfXX7nS+ff/cwmOrTAQ
9GqzXiuPHx9+6no/wfKCR17qegGZWyn95tN8gQrB3LQ10P+yZSMfX+x1DzwlhNNl
FJrPfvDev63EaLp1SYwGhrbBFpTkYjx+6Zf8bllHUR9GRe786jzNtZIU7GZ+uVA/
af33XFqjWe61gUVybQMUrBONlEw1vt6gxc5vIeeW3TRiXlWC2Z8bb04YlkzGw/wV
Q4FBMF3qyA8HROm+mre8+NYlugY607fTutpIO2uJphzbKK482vJAtuqly8SJJoe+
kv37ljEUk/FbxnExdhNykwlOMZFisnFYbm9tKwWxdP7taKzIwx72tRwfRxjs32Y9
7ulC2/KFstZhY99VxclkVLMf62zzVRxWe1f33sthVinNX+3a2rXciyZUNT8bYhyD
beaD00s5akAciMDz5AjjMVXGNuTG3tl7peueE8u7Nu5DJTJShSR7KSi8JQjSMKRe
Hcr8GY5KZ88K/VJkTZBbtIsVZlvDnLuPjD7vnwGJRzek/FQ/KVyDcW9eNzJjyDv0
vijPGtgtj0YEf/d7C4YnUK01zDiALQmTvQIQY+6oc3qLjkTMF1rhMm3aYy2+u6Qv
rM+zr7NkJe7OhlnbqkYnfb/58bzNZl80icR7gw2BwGQiplFOmgQxqQDo8EHJ+5PF
nQTh5bxRxg8P95j9gkoD1jQJDL+/0Rp0Ypaebmbyh/+ucQtgph6R36axiVrDj8ul
x5Oj/nsovOoGWl3JFyE8BOk9KUAzpT1PVozHw+wI3NUD3K32UWU2plAIigaiPP8v
54g6ziieXwoitRl+8lX6z1CazgoiBzfOz4t87FxtvDuOt40/iQMkhL4ljuoj/Kcr
2RRFS/0cMKS4H6VxqZtzGDXUESNbudjilyYazXNddvvGN8/AsiWKCUFsKiSlG7LM
+N1eNaldSx+ASRL4+FGYOAqHh+BRlOf/RWeUgUkILuNSBAydpG8uC7n/IR0utouw
t4LLwwy7iX9NAEaGxlfReNmKXxHPrAejlvF1EXYs7oD0kVM3HvZmGrxTCY+JS+5Z
8jSF9Ms2gpWK9PnMXT7VPeC5kuuO8wTVR/7mEXwm474ZhXL0oC1HGhen6x7zfUBe
y5TGiW1/poIpWOGb3WHBnhAF4Yp0DaLMccSOG/FFkHINE1O2vB6QrvAmHW6uATjd
R7sV9DQNxh0byZR8buHrzQ==
`protect end_protected