`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36704 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
DcaI24013a1ntsbbicG8fydv0mr/VV+pwsE9akW9oRc0pkuUqKIJQoGkSA8L8Y8Q
1HSM8SKqcTOJX3bN2tz/h/8L+4Y7zN1hv6yKO1zAFFggMcaEEvmaNLBK9FgoN+Wc
ygfgSJQnSEbJ3IahQJy5HM2U1STdyv95a6MB1Ju3v7xHehTOYNsqyp6UjTzQUGzb
RR4pSH+sFW4ul/4LmNdJ5JPbNsTXSrKTs7oZFzZ6R8KTb4gXxO+wtFRMcc1krkpr
fup1VJwyrqNDn9Lmu694lwJo4YM1lycCV0eaixvsPOlNywGURDHK0n/xLQwRSul+
kkX+u26U64R3XPLATGoY/kW3Q8C30C67UJjyx3ZE6N4pMl/ynLFIT47kV3EyX4VO
nElpXhB5fN3OyqjhRhApHoNTLmcXw9HUI5uU4LEJDfcOa2k6ZkylLcopCKOpc/2e
iScVGtiDW/fSdklGHNkznC6OmNTuYP3/mSRT8G20iUVXnyaco3dyBZdArPP5ehAx
a0jyDtOW2BrixFcBqTTo3IwUu3XFucdGw0WBV9y4xel/lWPsHAf78MpzhE3w0mgG
pubJKjupFFmSaME+p74m0xtbVLFn/ki+Ix9U07s5Z80VcevSBlhozHl3HV+njzGN
BAfObg7TjkkkCcsVyAkZiXrJLMM1hmcO++CxLVGnDeYp3QtKAbVlO3/OeJy+l1TR
gPZkrChLMsbZGcp8azsgxsWGrCOfGT7HDMCf+aASRlWhn/PbHPjRdjZtW2ncEgOt
qwoIJ0q871SzsdIjFb1MSZheO2tmv/92X1mRfl1kK12dTnyANYVy9dPmeFN7cHEr
tJj/oGwWq2If84vh6OAnsHYJVrEawMVpcR1TK82XRmAMb7REzQSZBLlQi2WQv4Rj
cJodBUGnJJz3IJ05MeoC9EDHiMKnASFEqY9/ITalMcVHmwarEElTos07r386OJeQ
l/FsxP+CD+TVgLru4i/EYnqxlxCQHsfLjwIxJab0Xhkbva2FuEhIJAy77319LCsQ
J2Y2Mf0qHqGAYZ/XqDlkuUP9vHGeQu4Z7oROeGnfdgQq5/7duZuEuAZyW0qgExyQ
6R23MuNA0jB7Jh4I8bCVGs7NLZk1dDTFTvTbYrA78LYGZhs094jqhCUIJftzTGji
0EFbPu22t3NTshcYBsPi8hX0DGPemaA/slsvEW9cGVadGCqFZGL6d41OUxJlcl1E
HC0cV2vKwMH5uetKVFbNPcLcObw7Jo6xIwcLEHm6DUcgWAZdq2MjmL2psXyMIdYC
SVLE5vXNbiOJqG0U4QtdJW3pW+HNp1GV0KNqisFfk522ctBLhMvQ3ZlcDQiS6FJa
Tdkv3JEJZq91aBtg1RE6+iz2sKsk2OynGg68YvQkubIN7LCw6+QRw0Q8zDrbiGVx
itGfbpYS55Wk/vAMUmQ8i+PAVdWXtoeud1Q/6TmYuDiE8/8MMM4WQan6ocQHJpwF
QiAb7oJFkddxD0Xg+GkXfGCSRbLWZNKIAAxFliUdsiF+MfbdgeE3vAb2eLkpeM2D
McjOyO++OeaSkMSnt8zxXnwUDS0vFSFZzlKnB+kFNz6NNzZCk0q2J2J6qQH9Ol4l
JQ0TquA8MZTPWeBiltJTozBzBtG7KJsGuyxCAB3qEXu/p9B75ysPUYuqswZrX0wO
BAlHifjF7fS9tA7tDg72ZoYAK2uIgD2FPjlGbYkTyAB/w6C6ky8Ac6tIXMdLO3MF
flZZpV8lC2Jyt6XIfs5NbyWzpW9Ar6jqjlQ+Qmw6HVbL2rJFRchf4BeoAPaNw8kN
0iZsv5bq9PbPmdxsx28s4VuJHsFW4T/xdc53wD/cl7rAHw9ATAO516PvuVd+J7wJ
JbPWEdoPvnxRibKaXY8B5mPPpvmYBX8ktnosQUNYehgztUEVJW4BQKJS/ghtOpkk
0ZWY89cpcq1yFYMuylzvyB0Igus4Xy2HytiEt38H1ph4dupmKFFX5m+yB1L55qKP
sCeuDJh72HDbcN6WA1WUuKBzhXE79igmUf9b/czh9/cYqJD8WJuVXeAe4Qdv1zfi
0rjUPb6Vtjx1foab6YLaKCf9/mtadpyM2+A5nvaxcLixttXZwsfZ9kKqOVTZv/CI
2kQknV6nchlCodIeAUSpWrY+xYaLj1deTtpxFfC1oFF2xI5fK/o3lRgCAV0bVFl8
k6Obnb3nddMq3HP/WM6CJDuN67g0GwZu3hQK63mTjEYka8v+ENzsVb3vTGayUInp
r+odRGFiYmyG8Cmzz0ci+TkQ+Yy77Pxnuma6gH88QOe3BuUMMUhVxG7Gfn+JEIUM
oaWFoNtFOC3JXD5hNPhmtczXNY/zhQfLqRiqDZmnM1FZsfB4PE0qX1eUcVWkJsyr
81TtNCTwmHJW3HQKTmXJ2pNIc+6Q3TuOyNB+yig44e7e/0HadiUk2U83NGbxbis/
uG+J52Qtc2MnCRcJOZAeVinnDM9IMX8d3zfskMV/V6C0uYey5qMJVHNSs9IHedxJ
SbOOzjrNeRx8QJjqbX63VjwEu42X6pqt7NxJPgHWDIBsmHvCZQUDKlRuJrJI9skb
sekL8PtypLbPvkM5PdvCYmhk2xOd/F/i+vIEVhAuHbxlV5kBiRc8gN78E1zJI8Aq
MsX0gPF6H2yQ5dOfyh+23hxoXtHgEYdcyFDeNxBHHSvwz3k3+Tw+MgF1ERruXLpS
UQ1gYs0wGBETh5dapZdTmNTDTbBY6Xe9OEmeXNF0a/GidbmxzBsOUPrqyArxFNYf
xuPfif8Q+7OlbyHDZcZ92FiZXDwZ2zBJ3EXYUOv8l120w0n7HZ58igP9+lUqi6/8
dJ9L41nTCB5R3r/N+EyPMYqBmN32jzEEksKl+x95ZAGnh4n3hY5mgxfupF6wW/FA
nyzUXG7k5GQKiztSpjoDFkPIcNKP4HMjrb+853eXlG29rlJytr0Cq19qIBiOMpYl
DwKuv3mYcF8wDve+xrQdEBUS4pTd7acSXI6tkHsUf9PCrb6/fGw5BbtU0pptlUIN
LIbohR1Gs6VoNaa5Oyz/yx4qf4hXqhGCsGyXEoVgnV9wXn67o6BHnjiDUVSuc7Kd
f2yWuI6n4bXeZfFwo+5F0/pj7BpNmhjhcjaw/zPs4BdPlpfoXe+NUuUhCznQGVt/
Lm1WJVDBk2ffF7m0LjsWhZCJWCfXIBDSYErHAV2mSnLN4ipSCXeAGbbHSODTRAJT
hEhPSMt8rzD92ZbBp71GmxF0bdpGIkjzh+jzrYYEUcAiHJSkNS0HOhAbSjmwfxTq
7LiqRblGGfHs0l64XY1Vqvimw678i9+BQQk197ux0Tdy2xEkQd/xEoK4n1ZKKvvW
N2GM11rrE6lMPNAyLaddesTmB245jT5zzdp0vevEu2f5HJvftKwukWfz7RVPWVJC
iGEAzBtrB0henzYXQhfgSPgXV3olY6o2RZ+vuRaExDxqefWKVCwfm07cbw4nPkE9
54HrQ5yB26tIqk9KKefh+8OkAui+pFTbJICQOTlFg3uGc6GfHurKoTNQX5AGULQ+
PJERtZ8XV4/fbi7U88+JEomuDl9fmFrOhYLLdM4pW5ERBW+ZG5yMxFM0hTYRnlF7
D5iGQiCTC9HxENTViXFnBy9yG1nZn3p1y5FcNIpvxDXL+mOA6Ggw4tokvxETWJTP
xDbx9Lsx8U9vfMR5ZR1n0h9vn5pUdwTdh6r+hb6pTOMv/HgpAMJITxO/WJNIl7FN
+U19V6o9/sKK9/ybzqHZXU5wRoSf90DLH+vnOXtxwFmObX4yJ/zJisYe56mU7Dbd
A4qjW3+/8vUiaRVF1o5q5Gn/F1oLKBY3Ym1RFlL78BnyMYuecpzVo0te83FPgarI
0CqUM57pfV+7uppsNhOPkBfXa2rWAa4stlxhhOgv5UkSdvUjtIF/OW9h6+41zw3g
Dk8DZzxIlS+DltVXeODJ07iLhSmlOS4GNO1naK3/y757bQXql7ddwmci8h3LcIIb
MG7VYVyznr/0iFm6eKF2eLcmiPMUyDqvqUyYDxekKirTqWctipBFuXGOG86ERDlk
+WI7Ce1f0c7hdRY8HWvYUc/tTE8YTtWWP9+sRQad+giJktSQWRuNJst6BVInL0zW
5tH5NUAwz4XBeM2sRTdtXXqclf/JoeMS6aLlggojZAjdWZGOkq8Nj1/l2+dWb0m+
Pjz1WBkewACHL1oi/0aqatXOQw/FVVAJJ1NjsvKQkXWMA4tf/m/094UuhNoSr9QN
w0fExOqb+T4jliA4TeGO2hh/Z/eCWLpfZ8iPDkP36bUkyyDrGYpbjiz6tS6eDE73
3zllZQw/r+URq6ASai1Cx4MPI6QQnCl3cntEzUVm7byPlOo0L6f/VNmjnCiMFIxI
aAwaoY1JqE4r+0O/UqEGnasWmCahuMsxVxVBQJDCrAuuGk212eQNxbZ6T/TlVK1L
gisBp6OYrPlDlRBlr9QF7JBSeFYNntzMU7I5+1HcTVA0eThzWWHaZcpux7PA9MzE
13nRcE2tnJtzgGeEPDHY4xOwmjOTK/cs5ZeGnSxASs0pVVdd2doJF/uDxIlPYdZ1
6UJRgYbjXilDHMjeCovPSH0ARislZvACX3TEneB3iA8am/fHRIXlrZ3EJ/2GvV/g
uLP3zrE5zEvPkDcYZlFoopugOhw56qpkdzJFsx0PlEmtX93zqgvY+Ak7XOUIn6Lh
pu6oCYh7MXCHjYbPsu9VfdRLjuQ5jSlJtNThDhB+vcfBUT75VCRJj6wVCP4qxTZ+
hAaWv5SI8MxzH+4ToUW77/8DNMeOxgIo26egU2cbOJLHJb3JGhH/025+N8wQF0UC
61rJy8gFz6mAt7fs4VN4xsZjW57+0zSkEMEmuW6j6vC7/ttj2VbpAPMOCUCN6rjq
4bzBdI+byxFk01YPRhOvn/zO0SYLw64IIqgFJ/eH1u14lAc+Tphn5hfcLwMYE9YY
Yla1UBEwHkzC/PflQXMTEvUpePc7QXyjy2I00XCASDK+YoK0bBVkGKGVyE9VS0Dz
/lAp58FJBhBetOtSnyTUEOkTSibTRS97MyBjhDoYqZr914oz+vhvVXhwmmmUy7iS
kklTKBG8rgqtJTSCnu2l6cfu7g3e6VfoPvOQVMpD0A7hhTCe/IZOt6gsxWZoeQ9v
pD731hy4w6bLzHjdWpXNyqx5u6buDKGr8CSqJaGzbXPC9i2w/gVdR1bsIqokZQHF
0M/e+i80BLr0wenLfnWhYnd49B1MuxLubs5A6dn22WfzeztyfdvZTSgYZPaFdg41
r9Yd/XmpU29SdOgc+C2wnEOVVylkIwJUVfX43TaaC0gYHsGmcl4J5M9dE+ZBHvfN
F3buMiawxPBbRY0yyvQc3Enx3lQHN/iATSIX2MwMDUICRtmTaa5rCR4TDFFUwmHG
Q4deM8unpfZBr+3N5VTK3tcO/jN/n8KeHxKmOFsOrKiCdKgcP4cUeh6yd0EPZpJR
/LassOeeW1CuJHmmGUzT3faY+DEp0IYUu3GnNSqauuyyQBlRzx/4Z3O0+vwg2fAz
zseDz8ya/ZZoQaTt6SAhNASOWyl59VeowP9ONLm5gDY7J13y7Qilw/nE5g2mHPUm
TuIydblXNJT4vfrtawPyka7srqTMCtOdaaX/aPlOWpKSjE5UOpJZkhEYmgJposPq
FqU5BTAPHZI0NXn5xuNC57cZ5YtLuqfVoq43sHvncBDR7lMFOebERzz7HD/ZtB9B
+RzZtFyuCuzLgeSrHE1MIG34SyGxvPh5pMoThdgYya2k62IE4zzn8ewCvTi5ShcD
1b7VR+jNSreVEYSJdmGJbSjmIU8PpMPN/H/OBZB/GZSxwTFTKGyl0umNRlnaPGrj
VeL5pfFk6fh2UtA22kU19pdpCHDeg/W1oC67E7LLHqnoJ0CEunsy9t+UE0d1i55Y
eFDywAPzrz6/uIp505eLoAgvXDx4M4/jSPdio6fSqfu/bwbdrtcj1pmJbiDrjAju
2Xh914h5/+lm3QETctAo3EXtNHQSBdbNOvzoAFkV0j3Ak/efFTz8Yt9kMN/ycF+o
gKr0Sm6WDKadlHBOiirRwNiRxqmot0pp1G6qONsAWNhh4+UK1nozQbzFR71xxfwH
6BzTKvGbZTip2SaxqdONiEI+uXxbrxkZgel80CSUDw+TeYw54dnDEhnJqsabn4RI
HkjhjfTetyXtOK21KqYlouyQNDK7ITElGFgFz+eTrS9WmV2qPeUST+pK1yEk8SRn
+G8NjxisfiZdEDtUppSBvUoMBJ2l6sCnKmh3N3J4ugmIY+fN/0ztsgCPypQeX2bE
Tmh8MgazVuG2k54tFIzkPXEceOrTE5BxBp7g/4J74YK9EEZbUoqqDPgXkGJYVZng
XICrJS6yoj25GRfNZDHUeH+n3coGq+DSjDzFK4/MU6G1hfYcYo2ozSVstFdZdiRQ
bCGawcMwa4dbMQuDpSz7Xduar+77nVbDX7xK0bBkmvas3mUdIJKTJRT+YrjOPVtj
XIFwvUqwSW5W7Fmm8EXmthottEGjZpMR43ytkVy2KdlaqBDnB5MPwlzi1tCngM8h
iKkLHtRcDSMk89u2Tem1vN8FT0Vwz22GKh+0LL2XuM2CU5EAqXebrVLogIaO2Bqx
KIaOEQn0w6P7wbEcGMnjOvVcNYrPCB4nd08sxtKatGpkhbwAXqVEH6ObxjOhoz1O
/DD9FII12te9s+XYgg2aja3QY8vz6MC16XDJvMWj3pSlmOp4CsHh6xtjQhbsFRnG
3h++QDbC4By6g4xYN0i/mdl01UefOqAy0bTwruu1okcyHU6Z6+eETul9O62yxSp/
GaNsPygREDYpEVaZZmQUBdz+bW1eXcEIpqo2S9MvfhGyuemDlw5ZIyUJrFBaWr8G
EHi5Auu/L7fFKqlKaghsvZ7Ww2MioCLG9xKl4yuOny3hntz/4iaiocqA1Ku4KKed
CPAHLnKL1hxyRaVA9gygTXSZhheLmI9PB7TFF0fR3yfKzMBysigXhE4y0SDKuKQw
SZEmRK7bhF8s7VACeG6gGvlazGvRhdmhT4/NlqlKVNWGeA5y3lM06HXCAnfcnCvt
iBtN9DJ9HhJTO8/y0QjipwAVKqXRvjf9qSgL5Jznb8bQk8fJxZ6HLQwDDlPozm0G
9Csw2lhp76QjfFrPZQ9vZULIJ2EQ4dTGo6Pcc6tdN5nBaifTVvmwjs5OW914w4mX
uxohdmK+BfeQBHzcP3JPmlhUb0qGTsnNu9KEZAxU7w1RE9Jy06xP3/WUqxQywLkI
Jg3O00sFKSjDZb2trMh6wZ2I4EFUCqGAPbPNZ/8Xj1hWcpSqWrG/FiEZbpaqkwHB
tdJyn0LPPgvljEGznlRbu+Cn97Z4gKyPr66Q8dJ9Ki6uLChy+DT1dgWtsp8f7nqF
z8uIYEQHMZ03G0dwChZiMf319vz0Grhnud5dbaALhVU74tyVAtlguMDTYh/eekit
xgOhTIuFwxzoLTwYBDVyP7cXWJUm/jY+W7imZuBJH0D+3FcuUONt2uU3mE3R7P9k
29umDfPAj2kiw65MVrq1wdigSPb/Bv4mlbqr87GS/6R3A8qsGFbwRX/Q2LKTX/HU
Ff1cJto4yYUauKw4oVtsb6xTEfIw/oIgk0FBFMxe14yATEmKY5nRfSSavqB45Vsa
hWCM+rRJsnJdNzPBRFL0VJgQBUoHAWVWzIqwbj7qrFUYBVQPCnv29GRMtK+MkYvR
K7DjTnoOD/j53kB/bLVQVMtZB3awFU4L2DFHNZTq5Z2TflhdbsFcofGUmH/DaHVq
kqJ3elA8HkS957aVcOycWTrFENAyzMszsqWx11mJPnc37m2GABpBHpSi+/Qgehde
V4Hocpragd+k7lRnho2cD4/gDaYG92poxVtgH3h8DSQ30BzzRTtBt+Q6fmQjDxvQ
Q0T6dt+cz1xm5fWOKMpxYJXjf98kw4qoeqIhL6lx7Nolr1sl7tZ4I1XJovLrr564
MoXEs9YIo3mTyAxl1DskyBBfsuy6mZ+w8N5rHlSIP0pivw73ygzWszYOPuT2usug
eGLKFdbjhG49c6K/gdxa10qBw8S/A1Ed556JMhkJ7lnqeNgRp7uXL5Ibpv/iVNth
7klEvCBVYN2/tAu6LthM6aN4ItT54Imf5dqgFv0sfi8OdVMqUJw492BEvmWUmnj4
z182pRlSP6WREZflPJRmi1KpKYgqNHfrfm/t7Q0+OKMJBTCJXa7zQzGLUlvyAlNJ
UEfv3/w8XIVNwPnnj/VHJLrrRgDNVYiPv20yusQ4xa+ljdFZkTt5yBjh6AyaxDWN
haX8Xb5Y9ZDu9iUUXnB0uRd0Ty5x77tljHvbBvuGdyuXeSojECIgO6pCyLUcBxTq
n5qWIsBSNvIdgO5RJ8TBTfq/n2B+EWy9DVoKBak6gIY/qdTTTwyzI2SLufLowB3b
I5fsY/mc7TQ7w8dsdKTyEr6aUsC3U9AoKc068a3a9+VHqk0hSVk0yhhlR7POCAno
1BsD92SF/MfeuTag+ZHdy8mT1IwEKbOHVBT32AJXd2DZKTM94ETvw3dn6pNnpoIi
5gmc9oaJthRADTUDr1kZRa1v1osSsA3zOYVdmL+eONVzotJ24XLKrZ59ErtnbN5G
e0rzM3afaNAe11PhQnOsvXSCvWHGvEhSpy+BIhRkWNKdA4LE7OM6Y6Y1M4oPkKuy
7c5ljBxSq69J+Q+lKiD6KioClnxXRxtjgar8ouhLd8/+xf1+ubA6XcO9gr3ypTib
aTjx4GZ0NunnJqNmFc9Re2GNTDxcOttiE20RPO/D0AO/lc+yCM9R6eC3TJGA3yDf
4WNJ4pnpzehy6tGXgdkBFWc6XIM7M67fBOdUwx5ogNMgi+pRheye2n2qukcZHt1P
Qw9s+L1XcvTwcq5lA8KOo7ByS8Mxyf9Zp9+KeOIgrbDGIjsLYRzetACfZMG6oL7f
zKjG5m3fkFUgpFHIQi5kjU4i4QhwapPfdsM0yftUcD5M9zgrv3FWQ/eZboN47jJo
0B6UaEii4eIITfVT6Gh1bnKfsNFToUu61ZtArbBwkPXVsLoAgBcG7gcdni72Pm6n
RbihXEwYL7rw7LZK9ipcAvYZuX97jl4SjRPY6Z6ZHbsXAOyjsrfRsIxsgMvq+ng1
6f2733rvYBTgTG3NDVCCP1uD6HBezrD2lhR7PN/AiRgNgN8Y922WUrss4z0qq8zu
eeJDTI6yAoFzxChUDuxAWMQxmbnxc4NMttDdUhBmoWb0zc5fr54owDeCKwdbuxIN
u9MNta1pbu3iyF6DE8MPQSBKLjR+HVRkPkVtH6NpGBelExLlIl71sLP+CwyK8rZ3
P52eMoNJv07qCYCxOyklaU62G5wZx0I1oryim4ijgNxIKhbypNM1HPTTTRaRi/Xd
oyKepPazUoP8ny/0kPoFED4sM8Paxw93MFhA+RFaZKHVpe724mjht3yI6w4UTENU
4k5ykyusfDb631grri+K933v+B/uKi3vrXF56qKxyLXG0GS5jjK4ANX3JVlJx8Sv
XZDDqM2i46+hR8XV7SfbmDIPgaKTYbkAUavZbhXpGT+H5dkuTP00NPElD9wOfyR1
rVoUjpJl5zBHXTU7bg0nMJcRSi5h2+xIKQuSWuV1RErPqbLr3VNJrPF16+OkuljI
VzY2iLz+Jz+8ssuZ54pnWHGfT4OJ69DLA0ibyNyhTrcVaEyO1Udg0YHWZPTIJjzn
+THJRnlqHN6m7LcrEoS/jfavpIVhxLBlfhfe846Lbr+kghWQp2ZhqTzLGZSkrG4r
nyJ4qarkXNG6nWkq9xBVgAhrhr/ftEdW1PvjnXUkv7HKzcXazXP4Y1LR8/rd2uN/
pk1RgVnFx7tvmBiBp4ADuxMHup/X0CYyayw4mby/9w4qFR315Jyvsmc8zE9r4tR7
Pd7e7gXCoHy1oC08EiGb0nQrjxCZiAXUuYiExqLQhqEnrhUF11VJhti97Ph0zyRn
pR9uMJhfTLfyNFWjSHWaaJ51khhFIgnD0lNdN90Xg3WHpXt3aeyc0n0pucYC+C/k
nqP22cWO8JV4xXe/7SRwUl/XBbEjUoXNYY0DnMHwELBoIUXvSVhFdLy/T/Cz03eP
SQzyoPuctRyjqSZFexvRgUo/2l7ugfbdON4bzyEzp8C3WEy/cFmO2BGhsmA8M0FE
bG1d8FDh+b4jNGPdR+/Ejb+42YRCR/N8/OMWxxmB+IqbIn4SwBJSm2+LSCfo7VaC
hPmyvIBdNklzdBiCgD11ii0KXgVV+b/LKECpv5TYzOh9WJ6eVKz46sBL3a7Eybjd
qNHllZPpWBZUVmRj1xdwhqc5QMtzUIr6qEnWI6kI8HgMoUAWMUrbvtAXy/34T42o
HyN8swX1f6aZu5tk+tskdd1HOeflIRT4+3cy2mAcwB2bXzKbYBolhXJ+wktm3SXa
H+qd4lkYgkXWUiDDxkYk4Gy0xQBtNbDOUfkPJqBUTkBSFwKksqOobXz08AygzZ32
1uzbaE5qNQtUOxgMtzwBmZYJVeJqBwckOJpYVcWOCcfs3kPeMU+Z+mTBXtn4rIXU
pIkYvo21+78tcPsUq5WxSB9lzIqLTvtm6RdnbUlimO/pSa7qjMGRBVPABiskkkMT
Ak+Mvdd9BJo13wUN3ug+BLKYNS31vtFoZfwYIYd2/spHsd8yJuqeLyYifFNeNVAK
NQfNbBH+EiMrDKGCQClByLJmFY0UZSLh3krMdv1CInIulyqNTJez04Q6mWSEY08Y
pexasHLtiqmutOYQXK0DPAvKXH1Rh+AxycVVhprDX6HrH3VWfuny0PIEOe2Qp4SI
B5LlvxeMBIHX3iGL1tCnvDW+KXm05uIOFEdJ1aJhsMSM3UMotTXxPJ17KgKEAVej
JoWIbKdei/Lo2QWi/NKS1jZGjIKB3Mh11veXFPb7u5M4UtIcvnJdnNdEkWoWU69Z
HlekBxPsQCS7uq2qEmFTbb9YOaP78Ry3f2VD2DG2qYqZbU1t0nfB/FATQ/rSCxsm
0yfeKshTbye2QV1ehZncrqxaEMKpDwQA59V07jYB9HGNY6I/wb9XfGkljYbqk4sM
52XnFR7NYl7UOEQIILkT/Z1AV/usR2gWb259m//Zq6tMR7nngs5UH4xBbYqQkmCe
vI3yDQ+bApGeWQqliX8rgVkbqDvWd7Jk20gqrUP+XIRrOsc/8Oy7XsRavCRKfIHC
mlyj3GFygKLs1vkTKaLx5fX/0gcAgDML4gDRbDMV4z6GeQO8zDXvf88cRmgJw4Lr
tjd5qRljlf6lrrgyARNawMDD3FeH1p3EJgFZ2EEIHkSTxC6lkPRW1mkJU8btA1Sl
rmzUPIjKrrieUJtC/1oDqE3zK5PQ2RD7tfoyx3pFAcSaRiAroLV1HkZ1BIrSVvzM
e+qDS/j3nQbb7T6iho5x+KR9lPbjOJvflOx3NHGQFNa6knRZEDnyciXldYU9ldXJ
x8uQjgOdQ2YFBS1CAYr5xMa8ksKFEPCa0Sd3UlXNq0OCwTGwb0VQ1d/0rS/+pZcY
md9LRgFY4wo41BRyaadIxgkR2rBLwyU4EKO+Zg33D3TK+w9CpWDdYmF4TFN8jKfA
1lyhi/xV8cM/tVuwF5cLvf4RCv6whMLfAw8Pva7f9MDRuoTDQWB3UNSAQbIwov3U
pVUrIKhA/kjpffR26nBq7mcGOhCoBkb5ARv1fYCQ04pXVMPHz/UlyVhY1wzABigI
Bgp1ZH2cPNRxTYKmadJqWMcgvfy3aooyTIji0noVPDHMFv4fHedMydj6LAnfWq2w
rjksUub2lB7BD6olfPUQSg3DQFewRF+pX/GPuDWB8EZHFqLQUfK2hRxTLGicbFUE
DNKVycndCi4qFDs/l4xWL2lcwGwMjH0jIYselJ2lOV1fu/3DZg74SFACUGzJgZwv
pZK7+/VmyDydj3MkYMZTqoUh5YoTgpS2eLUfsynQAR4IBdlnFf/RNSxSvzXgyTFQ
3hUDOdH193PFiRkFAE3FDv4GUPRcPoXOUaQ3tZd2+oncekm5R6KrgSdFYFQZq8wl
+0ugLZluQbU60xKzmNP2VXF+V20JJgP90u+3TGXNOCDEFOd9zpljEELs3nIYK/z8
n+314U4LL/ofKROB7QNCxBf+Twg71hY2jY8rmRYRy3KWfiq1XnBAlVrIRYZxS292
i75NSzP2W1H/yxr2TcLGehbLy7MlWr3BXrBoUTlQJAJ2b31drdKtfMKM9ecbGLfs
UKi2qqZa4ZMMR+2nUxoxc86DTnVpdPIu9IZ2TfePNDq2D+Wma4eFMmk+YD5lvtGo
XirLr9aLZ4MliXq2sJilsWEUVjEM5CFt7hPjSIWcGg3puNISG3v+wuErUTajjP/I
D2FtkPBQo1WMvfKG486N2KVJvYmePPISudHt1wmNXvBd7kSfBb+rqtfGhsWGt2LX
m2Grgoe7gaSWoT5S6u/4gaj5xF+xHFpecIf38b9aSa+mPegfwhC5HETEBmmJ5P3g
1Y1EmgMjDW53zuQEBTXWHsF9/R1x/XXJINjYMRjj2wJ0u4E1LgTB5rqidUoBJ5qO
6SAFNwb178UJSdjin7CZXWgdvrFW2Pxx1gogXNlfS8SZavTkMimbhudH6ORLU3Fe
EMKRDM1TpruflHGZTfb5SqPNY9B0yEtjarjPOGn+Is2qaiwphZWvSId307iPNggf
U13ndU6FjNJevpuCPP0i8eOrUepIzFTQ19TsaQTxioIIER2b+pPlC0O7BHjtv1xo
blEzu2b/ILnN8vEtRKwFBCmn0htXX4+2Dk74uR1LZiC1NX6n97YPQHMdvlkz2aWB
B0p6dSsm6rUzh4/ZM/qmaUciopJrhJUxtfg7EF9GyggOfjWSAhQhGml0Rngmhzbl
q4+XKAzgNPDnCT3UbUn/g5qCLwgzUjM+btQ7p7b8LX4E0mMS7bUgwPxmzCRuooMO
XoNiHexg6FqwZJ+nr6OwN0nEfgmyUPVhN3Blfxv97GgvsHoO/LWX4EXLTbv9YVKh
0SKA4K6Xs1XrDWZ2Kd6tCYM+eS87VE/+BLtMqV1GOPVu/rAQKt78+gIRR7DJglgh
vQm2mxOE3nMvcYD6v50b91+Tz79tuPsXk33Anl2XiKj5Zxkwb+YX1kPz3ZUsEcaP
LZkpzTP5ns8v+gmM8hbL0Ar59TY2x8Yzrg+NI/00DQO0vUdBxCiw0jW1cy30lUQz
zldxhuhMJxWcuCVXWGQIw6KPlpsSO2YKCipAl23JJ4wdrkb77VfgLa4qgbIg3ssG
FI1PCMENx9Patf6c6ndCMpNCPCPVeXhWIi5kQ2Cx1TUlqZkEV3RG/W/Ba2QGFCsJ
E369e0uVeqbZ6P3HT2RLx0q2nPyug/ar1w+3L3v1YtN8T1aqqOZa9QrlLG4KOkYv
oQe1n0AYu5othkuza5ATS5+0qwFj/7FSDf1YTJCZk87kZtqetnTG6YCf+tX6qLbD
sYSa4HKj1iS2S4+J58tedhrRwi33+lGdHxIQwXG7mm8G0VIKh89rM8VSuLYzsng/
ceIVRwNj7eAF/iwhcqgKw/0j+UJNO4XLjje8o51ih+/HKyJkqv+STpMn5kyuCsP6
WQ/XfjI7zkUgykDmfCV2amL1n+MWhGZuKl5J8d5ihZRv4FhK6JgPCMYIqzTAzat5
+eAD5x52R3npdMCWim/jINWP2/7BrkU+4TxPAnqz2Ne5+EooQNQ8fE9c7BC4OyCg
PKmzxJE9zlHDeA0JSJz9acgVPCYb489LpeiK/XutORzNBUvTiKQW13P94XZoO/n1
jXukGTQOM00/SQ/m9p9JehgELEQfpCD4LHjIz5Vd9MKdalkB40sPbID/JX8IYTM3
Pl0mcv+GQJFjZVrca3lrkEo+AYBQ4p1BFgArV3uiihV0rK7CEhfX1kVxEdrV65K4
b2+CylTVc+n+IREZQhmQAdG0uLYMeM0SR3GK2D49vdoRfdBU4g+JJ6sLex5UmnG5
3b8pnUvJ8C/SH3TfPUnvb3LV7FpkW35YocTE8f5PVktMNIwgYZoEgWAGD8hmrovd
qS7tMv2D5InsANX5128QoDrBcx+4sPkgT/6D8A8NNS73bndQp1JtHdeGPoQHzWxd
2hxqHtx7fWvQyFIepOnkgCUNgcJ4yeqQPFz5vPZPCD7OOuuO2vwUPC3I75lX/q4/
VppSTCZc5ERqATMTQzxs73j0CXe5s4qqIVDIPagkklBwQEn7nZ3+Sa2eMWHacyB7
UzDO/WUmadvzooika4S5GUvgUvljyMHtdC12n0D9pTxOkY7VtgQDEvV3T8YRQP83
hyEcYByziqXnLWM/lmouMTddJiIkmNuvtb4/mrAwrfmIDUEqyx3F20ALZjW8ffe/
+gzkvU2+pFh+7WdeDU1yR59LfL93cOa566LjR5KFMD+cJwcrJO50Ojgwyz7tGBil
iKKKK6ZLmcrNomq33gnA+apB/0YIjelpQibuuiOz4Y/0SifVUJAt0n4eNwZ5fAKR
kSQfKsU0L8HO7o7nQA/cZEt9BWGCNQvQcZPMFZDpZLG6Asm/mB56V1spv4N6kYOd
Vb3/l9UhKELg6Ma8ka5vUmP+X7dM3MqnazxZ3naR+2Qtoymo0+2XyH6OxfaqCh5B
ULpZEzkK0JXr+pPPk7xBDmo5bdPshgTBmKYauCdAYP/i48i245ernzMvC6iujjxe
4Hm4V9lCYvtj+quWY9RAHNNYdQv/1Raeof52SR3/Bu0kUUsW6lamW+cNeNO5BYG5
4/lDkK8Ko378ZVHA6sKoTpV3U3jGAOPnldx2fXAAxTEju+sbtIhiDBHel4oD7lOo
AKvyNNSDMye/b/scOKXjxX0l4phNa1NKMD7ARMVoAV+V37JyPr/XrwE70DuP04rz
DNuZY5vHXAmRSkd+5YqiCx5rEpC2BL6a9ZObbbIkdDOWZjPTwpS/vehgMoUemOnp
dj26KjkV5xofHaKwC7o8v5hef8kx35/gBKqzB5gxdCYZvHkCYwTAvOrU68dgezLH
BsrbuupW36uz/O9RfyrM8pMr4snLfdACNKq6Sq0WGLIVqbK3CXi7nwfeZ3RjZ/26
0rAEj0jxfDOSW81dcmrIHEidBD9+6K37zP0jXm0x3F+7jKKD3u7wevnBvJeAzsqd
pa7lj8YSX5Ftn2ajJ2OMllQfTTTBR59SNuqlnSR+siMwha4mK8P0vaEnFyirdjED
Ko98fFcYwVsmgrU/Sy7ORYJMDCG+DXOai4r7c4YbnwV7VInDMd1DQwHg9geLl5jm
IgtMX+gNEXAQbt8b7gX+DWmZZTz/2Ja97ISETpBIPP79vgg+kMlgLNakJhIcXYX4
Hkxjzhq3z+qB4l74XSVqQZgXIOsNJax8H6u4JM7J9fLJuNjmqVkK83rlGkltjgVb
OtcBNiUDL5qwEtoCJXMmKYIJ7eBHyJmDeRlKh63QAvuP93PWWWhzNQAFumgWXpZA
cPLCh69YvvFowwBfIKLf52yaY458jiXbVpniUMcGVPXMMWHOXZH7UoIaHMJzRdx7
NhiJLwNZOCKKFDOrqWtAkxelO4tjXlG3UjJWEN7l9/juJUQFM7iaiEsE4WaEj8RB
t03X6tsXzrqmdRPTbPNXYglSZ7QCfn8AiJ4roT/WENptgBSWZJlNAY+w9qjs/fjr
Sy1VF+thkxNdq5YotmecmlkUncR+lBhBo1ffJoo/gEh03QrNQp/iOcR1sDDFvE9/
fcEmiHX6RGAYX4JJbenZ0X8uZ8xuarzdRKHV2yyMafUnrFRs7VCi3fAUMbZYje7t
oKiBjB8dvCfPHfQhPFiWZpJ/eKZ+Ozv2M1Iwq+AzaijqVVgCVw/KXs57MmDsS2Qw
TeBkI2qdU0CDeCFZkKcH8NJ1h9LTHhmJ5WkXs/bUketNqRHqL2UiRJQ1eqTPrwoA
hX9r9u7CSz0W2FKhY4eOENdE8MZHNI82mP57OjT/dZ8xEjr5SjerCFtyEtxRo91S
W11ph8pGnoQzxVSDtTtO7XC7CW0EWU422NLOCJKcne44dwFb6Q/8J7tCuZMO8gxi
TIsnp116Vb/gYU5u0PyWTAfiAklmSWWRgL3zx3tM6mt98I0K/LrU2u8VFCpvXOo3
E4hpkpVQVFB1srBjm5bxipcMEq3oXfeg8k9ab0IFHwH7RAFM81J3Qd9uzPFLr1QK
D4aft7TaNR/WlaCuzs2hKRk5enKhO5YDg1xhB41FNoj6eNbrBDg2FWKAxJKLsIjZ
UmA5ftq0gK364cGxjQEm8lrXrsBlIvF4dBVhbBQp+5i6z2kNPv3yiBkY13K7EGsE
C7z63Je8n9srZsiJIjKok3Y0yqupoVsKNyJRdronriuwH1sGMcxPBx+EcVhz38C/
ak2ET+vLxNSHc1epD+nxTUpLbAZTO//s+rpRpIBpm+k/a5micR2RXZhTIdmvVoXJ
joYVWDh/jJW84af3WUmJQbOndTd60Hmhu/LPtAlYYNLN2pAiJj/7+NwoNsU9nzX7
OB632FlNflxLa6guKuvVzbOBW+YACT1EOaO2xSeq0XRBwBu03Dej/r0+icxWiRPf
0tjT96jrcItT5qq7oOQYZazqR9+gui0tHN2tRWVCsU5Hw+C1E6yv6cXTsaxQtKc3
37QblxG94wuGKZXyh3l/rfi+rLWMayBliB6OPCsTxR0lWunc3ptFTyrRyoYHUFu8
jf/p6hu8XDNeGKtk8MEnTDZcGP23NcqCTAwRQXp3TozybgaCzY3n/m5Mkyo5aYZK
tSk0YjmwVfuZrEYaR0neBpiu9WmZrbJ5HG4QPS17KQhYwoeEBWWOIy7+uJF43GXE
1rHs2UEW54HDxQDdttecNx/CDrRVeJVT8k+urdQBvEMqdvO0nvYyHF2jHSbZbmFX
VXO26t9hn5Y0RBOc+ZCbh7mQk1ZQyI7XAW+PzqD0WtkDvXFXiNxCufylVUlJxrOZ
8I00G3gYkw88nnaK9HWXeFOypuYuy88VPNot6Rdhu16pydstUKz3Fx/JCTuIGEXw
U5x0lyn3COOzbMGGQUfchfLnRtjidkX2p+FSYwdz5mKwpyzhfIpmHhAdII8BUuOS
7eyaWu47Ph7iFCP1iKTMU5+7yNQIXEvPMrQyVUc4j8JusK7rygzZcTNx+Mx/HY8h
2xWfJwv05hQDN56lCYkAD++S/FjmqFhKfPzS2r4ngYMLOF2I3+zGrYar/j5XygZ3
0ZsOAe8GFzjEEDo8jothi0Y3UX9QkLCl9f52z9un2Tm5c+farASgOhfVTAtYNt8g
d1jAU6E49HgDoGKRZojUC/xF3aYbjNPxbh09Qp9zTBJQA7hqjAByn8HErrScvtOu
g8rutwQoztYZ4wWe2kYXtJvEAaHZHuBXjxt6vET3nMU8sIwA7QPzjJGXf789PU6W
+mTa+W4DM+9MPkhl86Td4d/iQqFDLzpgKOS6Zp9O6veFpebWc9FK2BQ9KeUU5EKI
ppMwCL60YC28dCpJxV8aevd5MD84F3Ij1Y3I+5vjvCv0MDqGhZc3h4cMEtgXBvLL
jQAleXC8hb4+LsF08a0Ed//W5/3UgRlb1JNB2YhjrBG0vPZnwADoCI/XZ32Ap5Mo
UcJ2SW9y7Kj1X6CJqebYR+t7wa8sp0nUXGyoW/l/+jFQFxWnhZy/vwaGE8OPy2w5
jjOvIB0HZz1/8anWeRCJeozRUGNNaY8KPAigvfWhaumDJnpZPF5Eyq5oT0OjEy79
Qqz54THZCWyPFtmHGXVv9nTQCJ4qAsCOo+r/DsV6Tx0rzeqv0aDfoQ5uDmjtm1VX
kA1imYQ+lORWgoFKNIn64rEaL37uzmy0AGyKrcsdRFb7QfQd5NJuo3TrPsKZOb/D
dHLCZXDGEvgO7FO1TX5IP+hNi5JoAbblbknu8mGjfMxnk/M0BI95qt3Z3SBPSqHF
ecRE7sG859Vfvi+AFq/TtXoGydXyMDXexkiyjKT5chexDO99trpEys9SeURiFFYE
0z6V3nAmNYM+Ar4y4+kGWLbaE9RAevKXsF1y58KxPNoMHh/jdlffqtuOROxE/Aym
33ceyDaca1rDrHRHJCcg3iS8CwNzJ+kVTs/T3TrZM8/ehUuNB7SCdVSzseLFb+hG
E8MA+9QDbIh5m9QomJY2YeThAQw/sTkOMNluaWaP9XnEH33joYuhz6aq50ppLu0U
YVUMHufyR0L1b+0Lr+Ap+FcJTMEM4uyUOEM2YMdEyi77b5Ua4uBU+z3+aRcKLbGx
ccm42HzMZsqklR+oQAt7ynG6PsgsNpcce8kxyoKNL5TUVByIScsq+SCpQuB0wchk
w86Jv7nhK7b1nQVGQABUN85V4I+IA4QNw/5mDGnDmXSeZLzA64SV1nsER9B3F0lA
5Y1VM4gZ1+PUKdJTKYtMtnzgIajPVVzwXJAdhRQk8b4+xtWDy0LpiylpIDiPLSZZ
4DCdfHBDaT2iFTnI32vUF6jDXGLTmI5mgZd9cTsxkwGAkhfhtEDtT9UEWQ8KjhiC
QC3c5KqwBJ7n+hF/v2JdEDE2t1/GYJAhm3snZQ3iiujtUx8Ak9DZlef7bZ6BPlvv
L405RNV6WsQxzu8w8hwUjfTtSqPbMGPCrNSN/8s0bS9b3sSQKBw5+MRlU08FfNK9
jyjPi5es6WXsD7uVLPoT5rhLDwqvu3Q490kk4Os2AR03sFX6ExCvS3yANIQ97EWi
vtGYzgiuecmA012XGKnwo33AEr17ZL/p76Jm5hZnv16JMlgNQtsAk9FIb/Cb/cPO
S5K8bRrg9QA/nZLZz8dfyTlVlLyeexn3WVyK1x1L20XtsOG+85IceReOxHU3O7Ti
S3Y3jnRF+VClVWhheCriYptb8+FPcypvf6RClf44y8/Zu5vuldMcmglLrRh7ual4
BNWC1SeSYGhZysX94I5Va2lrXhZlug4OxjYOEc1mh3hHrzmU9h+WP73F1lhbJ36M
nDrkANe1uiMNjKk2wTzyiiAPYHK//Ty8is3X4BCbbqCP06SPQ1yV7aVxDZTN7D97
uALCOg97/fAUgPcFmUFwfzxvTBC6a80YlPulal3daxMtu1aCmn/4MzzmOQne1hm1
IDn8Af3yRmY/DSAbmbkpbhGuICwHa2re3hKrC+XfGx3Fjm6Kd6hroQZrhfpYP8Mn
FX36wQhJxfys67yFUKlgV3TctKj5SYZae+0IpWdkt8bF+MEVi4++xzB2DQ3cUHkU
S4sBSTZ7vfxInQP+J6MogP5+PDUwsqZUf1+vz27I81ejZ9MmAfjO1BGI38tuIRTf
TeMOBPa3UcbSaBlrfLZLULS9HmDkViWSBq3OzBNXpycAMOeIYVJVcDJdPGNX/xYh
VGLWR41o5YSePbwllsWnDCd+C2R6hi29hMLqzU3zotZvZ3Mb0+tZKviDMJVuGN2K
waYZ7U+c8aNnvCdYsagnNnJCEy5BemsYLO1iNdehS1vPnBTYF0Hauzs2Hkrk0OTZ
mGY6AKLpqQuS6YECDWoB+dGoD4cCQhnT8uVxVmitdEcaOrbgoCdBfvspRVLyL5Te
CoxNLapAKlaz5oNNLnlInBy9+gNsEAih76JXfGvU+gzgTIjQ0u/3ofB9pVDgY/v/
Gz8Sn2/94rvNjtNiiT6laXlPMCvNuZyQGA9tlGMVPkaNh1HNLnwbLlp0jipoap8v
7CIHY4DCAbBdttf9XY0yG2nlxWX5kxKcNzO95PaBP7aBWRgaFcaExFgTWqFN6nl5
muIGd7duPNXYN9cF15gp+IkCi2cPAP8idDZm4IBL5FLg2ZRyLUcQ+Tp6zi4kzE+S
VLO0Tjiil5cFdXXcmr6qE9NDThFeKB4apC1Wu0Mh8vZTNx/h8f7I3GEKJyrVRfX5
91xgArMOvTO+sqese9M3ympXQaRpyMm985A9s5ZUlCAZvvq0GAwrsL0YZJt3DdGq
sS1kMrXGUYUbgaMcb4gigBrYYPd6Cx9row4+NaApajFbSyTItvW9H4FEZKE10ZMS
BE4MJMeyL9WpHR+mvp254a/xlkcpzFGxnE8MzZ2x0o2YsEXwS03frUAXqq9cz3uU
wOD1taWr9g+/Be2n579O8rfqJlVmVQj+D9bf3Lnwj6/lP1e2+Az8FisPK2/KMUCO
AsGnwZOC3vZRQo9/llqNEHbkVOvnopwpNJdI27hJb3HoJTEICgrkoQyJh1VtvoyY
UcW5Be2F11dSjAUJwkY92F01z4x4P5hUhuG9igLlARmucVsEDVIH4/H7IswhXBzE
KO0ieEIQUPVVa8cW6hap8necqyfbWbHayWH8gUgPdbotViWhJydhvYpIoHRXL2zO
B3gCHBXjfOSdoRQi1RDxi3mQdOAZZchhbrs2gzt7DZ8ChH6waI0BEZgocFbavuA7
u3hGjbbHIIbCRhLFZXivkL/c+at7yLkjXHjgIMtlPq7KHIT0MOMelkS0iMtIQksQ
VeHnCck2gYxKGak80WHMjDyWnsIBIwjB04d61HbXvTmAqezue+CvMbrVBKQafmUo
UswUTbsXiAJ4SVlELM/fj1dss6lQQ2mkG3OHZKL3USffmtZdr8o0owb62j1B4cfn
tC4T++U66z8eZKXDuY/oXudp60SVyspcxZuq44MXe4T1UOCN5GgcNaXSqEKv3khX
KTNhEZzhDFdEgS0/4vkqKqDdGZuZceZR0WlQxOcYBRFlPWsAGLM8uN1gB4GOoKYp
1EM0d+ZPv18fKRCAbDSJzuk/NpidaUf4g0mRoC9x8rMnI5ihIxX8TQcQdTXs7Fpk
vmJBsXTMMzpX2pntbw+RcBMu7SdABqicDRualUd9kkLRVGUB6xz8U48pCz0WHsnm
TJKHSNZ5cp9809kGp0gdNxhXgFejz3N6I9msvRehmA2S36WXhY03TxZVRZBIoaNE
E5Kq3YYRyzL61LHGAWsitXKsblh1ZNoVYW/AQajVhD6ppiSHaDYIP/PvrHBI65V2
2kIpTZGBfINh+FS/Y7UxAuG6cjE68IpM28i530P5x5lwitBTO2zZoKVyDct/sJkv
CFCC/VrJ2ErwcV0fWPKK1tlqRaf3TDKE+7U+ozqR+7LoN8eMJYlANYd7aIOnyOVn
Rk9lhtpa0hXXDn2HnHl4AL3gmvHdGBLsW3fp42B4kuekFe6HEdYMt4Ft60otU+LT
9+KWAaW0MSMLrK+VUwiGOQNvh2Rcus0AGF9VEYdway58zubv1e5U+ICZPeKN9m1n
cEVQeorknlaB5Ux4kcqMS5NprlYjxQ7da/Y/y1TTGFLCeBMIfavFH9fZ8MKFiNbg
py3DiyINwItg2zS33Cfh/mplPdiUQz5y2CQfdES+STX/YVrFbtjE0ZBehSFYG64L
mRqtqX+E6+v+f425jy/ymo6KfBxz/4FMowLKEKNPsh5NaB5l4afKChpbHJXPoUvm
nGPsEm7Gk+DglXMMKDhzv4UHH6TZ1rqhNxgNV72lAqhuAtNmhFnGbjVfaib5Rg77
EdQHGMbQisM5r9c+IZ1c2oMG0MhJIYIJouUnm9XhDUZFcQ2kkpsftigKj/fPMi6o
sE49/e4rd6wWiNhZfX/P/grXy8D+KlYRm4Osm8DhLbjDIz3RzYVQPW8M0gUw2Efx
CCi52jGcm8re6DwzviyChNG39QYlAx20yWEiusLA57RDjWrKlfs2eW/Xb47BGF5S
9YnnWsHp8j70SD9WS0AR6WJbkSpi6aIQX8ZAnxsApIQHlyxp0kJvfkB9/YEt6BBX
E1tn/btveeZrs/UQj4zf61MgW5auIAOhHnQUc6ZmX479w+n1LJ+nRUikxPIWO6aH
ka3Aq6tUp0vegTHlgJ4Jk8DUwsBIjPzpDkW5ejKjTLssr7BF4todM27d0Z9t73d7
kHbPmF37SdbnnxkLQNgmjd46YBE1KleIe2DasKY/bOMrzMIjJmsblJZMT/vd1c2Q
IlZYQy1vv5BQhC9JHQapLRDJgJ1bRNBXGM+3eAohFsdKCFCM6IDAnn3Z9PJ2lBmW
lzGPXuDh3QfieOKP7gUJtw0amSIUZPILzuWUEzoYTSGKwgsrYePRCMb3I1jcZEEW
gMTNI0eN42e6hjcqJEXTBTU/VfoL9up1Xr9TbJMBwda17xjLqAG4gHLMfz8aSzud
YFD2zmEqI8RMqkmTXKd/zwC2iSPhcTTCd/8j9aunzNhbN26JDclWQZeeFusEihpE
nL2e3pelDECK0YinM/aY/N6noF2O1vncYDeakdpJeslccaI+YPuC8eXQA/p/c3qP
nh8esfQqSjjZ52/ZE5xk0fXvLGZKR5/GYzWxe8BCK1ASvBEzR3OybKTuvwejsNfG
4hllTRQzCQE4HefoLaIWq8+V9sSo+UIII5CAOQCsekVPCUNh0P5EneKk9VVlB63Y
pIFrB6XIO8rdW7yPQYvValAB7wc9DQpfibInPVuZkrgJ1YlL+8yATVDBy+tzRjpQ
pRsz7m7+0+Gd70GvNoVPb9MlaTj+yjiNJu3BUorfZxRyvB9vR/sWjb4N9LBHpNDs
O9ZN431gViIqSBOlQWN2caL7FV4D6hQqq3UNBlzsoJCFs7pGwQAX2z1pYxpWTVMv
AbLaL3o7Y6ek5I46BwEL55aKk+DO/K7CzWpg+wbLqv5US7n6+5M3Qe7lrU4n/Pva
VtFgGjG73CAE3rD7TB7f7D9eKC4Kwsvqgkigc/YPXVjCQb7c9RQg2D9LiijVC/1W
T18cw4il6rU+F+gzEK9yZeQxuwtD/x4CmdG2Tb4X+44BZsxN8E0ao6MwS4NV189J
Kzts0i6bJx9kZgfKuUsreFK6lYNPL+vFl7jvKLc5ist3oEkKaA7iF1+a6NkdVmb9
OZ5ScnbcrZVB9WhuUgt2QQxBY+1hWG/dEc349Ez9I8tMs6r1De+U+wHy82lAcd4B
F6U2Rk2fedRSqyHV6G9KMXiJFi2bfqZz2xg49RzJGwWvagwF1BJq1uxh6mkE7L2Y
SuYSdt4KR2sLc0vTt5Es9z3EUtM6xAQYutXOYtAPIzIDY+QWP0tS1IuJ9OJQzSoV
gfm7ud0DXiStwkB0I9A+6kL/e2cNZqyODhknBE91jD7mlqJ7BKb7kyTMJ4mylQh4
Y5uH8rqoyC8YLC12EdWuFk3JocsIKbfSy9Y7Fz05ji8g8RM40bzFXY72oZPV2PCR
Iqxx11QniVE4ZFpo7HtwfNc3o78aNUuKeWGJxgHrOgyXp7Mek0AmR2tLBR+M7OIU
XcbixvO23CkBQLtAZPzattHLtgQUefHqriBZPYC8Qqkk7z9F9FcLdfR5/B74khmQ
vtEXNIEGEq4bL6B52uyOz5saY9SKjPhvGX8kFMCa5UOd2z4KBgS+bS8ma9zniGQg
YgZGn12KuQE7dfmzLYvjWoRADh8+UetNv71jBlHg8K29fZzLID9BFHo0tKXbT5T/
Ox3WwBza6T4d2WRbuugY4H3gxAxJ4jymsEkc5qYHk1XTJEzqalo2pYZ2ItpTugjm
6uQx4S/G4y1l7M83ioVuon5LLVnmV48U2QJ0yHpiS+goyR23v2tJc7K5XfcCMe1d
x2JAaevWdgIzUbWPYg3zyYKRLJX1P5F682Wmlim6SDr6oCUt7IxutqJeXmhrQRjr
6vGBbxnIoan9OOR7Ntp9QRzKLdPg4uykV49K4+uG4SbB6nGk4VngXWYdMa8brXdC
ymvOgrijXRWiI7azP6lm6UZA7zsdxhZfQFuU51yJyGazxwdX4r3AzvIFCiB2oQnr
41bGXqkkb6BxJ3jtRY4GbDKy6heFYBSalf3xb0PPu/RtDeUeftayq/ubnPpXPThp
KdXbMkcX2HBGQn83X4stGIwNAKu2uk+DsliGb4TXEwElwM9uSh7+x5lf78k8DTYt
Ol6X06bmNCAXvCnrbfAIVLwP3WelLgTY5nRaErZIe2/vd4f8yAHEoL4tiyDleMdH
hZvJLnkNQW6W7ljvI1sALdUW9DAysqpURcXAuhQfnJVWewTaejQdV7RCWurwHhkm
ji3tpzPPAS8WZ46reG57uSAp6FJy3dZYxFxdms0CRWwagR0e4zDzfdAgj9UGft2C
/sknq2NGJ8Jfmey3nN7KGi6+HE+fvzLaV5KHki7uSOVEbqpIiLsnv57wOXm1CbJe
7hS0BwiCFIfmlm95RYfosm23+d0MRuiKhx5DoVAalPYYHMLyPKxBU+/HcqHnS3Ax
0/262edyD85V3Gvu2dp0Ri+E+Cg2MKZHqhKXpxIo5Ht72DOs2gCOGwn7zuvrOXhO
L4y65rpgM0/Rav5+H4jC/ZfWIUiAgkoH+XwtrOREGCRPTWv2MHFzDp/zvrZ64Ac5
aKXYwEOI+agQ5EXR7zVJ0/TXYfXcLoIK2VxTYTV0C9NP+5cMd6Bze65xn+ut2tfc
Xg6wjaed7xMOAsF3V9LerEL3oIAw8fiqglfSh9YNzwq/QqXyFGXBSfIopP1/MWCR
XXdPVg5GMchSAGF/dXnyUR2uXU8gUwAw8pST3latvfCC6I31smYA8hpy8S057L0V
hzBGSPQncJACW5+L4uR8bOxuLnu9evDGzMSHbGXG0P6vr+FsgG5DGu4jgSVQ2lxd
3ASh4I7x9u3lm7N8Dh3qdPBCyqNuIHE3anTlGie3Psf1LRpI85NsQedDuV1HJO3w
2yhz0jYOoMR/tk/iWTcpJ8S/aovlAsvGKO9PeY+Z5ZAqf8p5AAEmsU4cTViUnIo7
YYSUmsvz3S7PB/GrzzGukuLeBt3yDOMSWQB5e3GahSIDzobR2nZij3YESVUfPrtm
9GNvZHSPddp6PPwppB74rIKdGdV9QIayZ/w2idXYk1+g+TbRPALAUH4i8E4QuNG/
LYiSa0MkRl/GhAE7VJ5NK7q3r6lmn+GRyhTwNFRExqVw2TdWgaIsS4LMPVV+Uuhu
aHtWteNr13k0G4Ur22tFifdkqFQmZ/l59eXmgACxJdp8L9iFe1FacXWGFLLB3wq5
VbucUzL45/GieeCD3wv7y2Yqb9nWa3iihu+mLs6KPfPyX1FjkkC41rZyLNWG9qQU
zlm0+LtJNrrZfMiJOu4zclUA+lWyrFJzQIHMUq3sXF87cyI0gE1xMbjlTJj3PhQM
10MS7K7uhoaAXBFfen68SiAhU3wY1jpzFidOBXxiU4Z4P42lD5Tkn28IIAzZL6+8
Qgo00TCwtteqoL548FvhU8H8t93/vlPgeFi7XzxmawWr+mgo5HdAziRAdRpumbcZ
wg/1trfwAVBFbciKvGyuyvVrT5CDyNTkA1RqdBY0Rp35Gl0Fs2oc5jsQLO4oLtzQ
wsoOlxx39l07bUj6sK0ncw2otEHYO4eLzMOKFNusBOy8Fyhqka45prptFIod1xur
RnuYk/OfwqF59RR9uecuGDA1nLOHoWWNZ4Gv4QthY48Ig5OZ3dH09cvpv4LDjd2v
sh5EeEirFAGAJU22wUc+sEOAce+6UoOwd+FAXTWkkj+xKyC/fhuU2gnc0gPTkFiD
1xUGv1TUhIeaeTwQwuoAuWTxm+9vipk6VAdb7KPmV4+igwntpqvU8bGarsA+Pfbw
I+4dl8pnPQz6Af3cmvVVlswIHUh7sf/nAbInFjjU+KGNeph+YAg2hp/c5aBx57+k
V6IuJMdKZSthIlkkkL1JEeJBO3dxkupp50vTgSI1YGg3lW9RnqlLHYPt3ygFx2Gw
KtPpAKbbErr7kdB/lXSODKRWmUeZqqC/Thqs8YnoAoSW/wIvlX3VbpVuWjlTeLfC
4PVRNzu/K0aHLN+MzVTysS0NW07m+bODo053A4qt59yCUkGMGXsStYm0Gobj3mUP
qxh6XGEc6wSXDfqxDIc9zwGMxVEuagvPjTcDlO+OoFoGdpTxmRxJeuHPPdpTCY2X
0SHaCp15J/vcXo9gwofDX+ZWiKLx8Tht6m30CdhGFi5KQDP55TRuQ41P1K6xA24O
W8LpoM/SSAfBCtFc8NuK1Ab3zt69FmuD1nffkOovXebQckUWYf77AA3WlVb4WFuF
CFp9WydHBVszh60xoaYZK7SyHYrK+MnEY/msdjVlT4Tx31wtzCmsz5KKuPWuGyRY
8+Kh8Uk7r5F6Iso2upaQ0knoetCF6Dqy1AhHBw3tV7W7llVkfVh/RdCwQZLj4TTE
q1y0Jjm4jaORAqisk1huNLuGFuhHFswAJl8wnEwzpM3TgdJbuTP+zedNh6xyELOo
oss/hc23KbX+Idn4YxjSB3/sF4iKEooQG2RmakKY8lCQvsJI06bA9YxwY0cfUA1x
1f/Yu8nSQUEpLciOcM3VVXUCFHvtmxHNGbPe4K0s2UCFoA5SOTzazB8Jh6WSol8i
FIhP9o+t/0BOkSO2JMqlWXX9Mo5ZrAo5+Iclvv8NKaian4OKz2q2AQaaS/PLdF80
ckZDhiiAskzNOzbTlgA/9+xbGnIEsu8C84DGeWjXiel8wPwzg9rqTQZqZWPx3lE7
EcQfoE6b9dkig9TAEB4UgpChRm7xyF3NUlmWAsZ333ej2Z1HME0FVnaJwY0l0RgL
eUXv9lA3Jh6UEZhq0Pd2lWRG1d4EL5Ge2U7D2bTnYvCEHqyqn0pteKXgC6tMGbx4
7f8NmmbWO/gipoTwRUHzXU46DcbfFBoHq9OpeEfxw98AJvOHcjzHxXHfoPqU1cHg
vNtFWjR7r0g5FJwq47CUtYPA4xhoc8Q8rE2qn8TFCsycwzTaCJXjOXP6vhqtNcwE
x1qPnOOv9zUvBO/KKdQ/18Gtpk1lPVn+NoXFAJ9G98X+xBIaLXbxKpa+Ay4JYt29
D3otN7Xn9pkRTEFLxPOyYQqWgwGzq1puhG6nfhu5uHSQWuyPpzKHJa2oljIb69tq
/1SkVae8UR24+HlwD0afLsFwN+FFmcnoC/XEtccMXopnNyL5BzWRrIQJv4+EEXgt
rbWgaVZfnBKpKegp3WnTGGwOTJX2B/zJkqtHu2NuNsbaFsLWNa7q6JnUIWEPU2Tf
WRoyh+AWRY3zuk+Dh9znZMLshL+UrCGTO+lXxviVrc6y2lcl7j0kDaQ9yCmATuGr
K1SQyJc3y3QRSFh70QsdIQ6YREejoFMWjiUxrZ1997w4qHpOKzA9Q8L0uYc7uNir
ukmFVUU/Z/JJhPgdiu+X/nWFpw9zBaEXH66Yw6168d1CjpxypKZmVLQYtI26Sgy7
n8GqIpXcjMPwMbM/PDo3hPOAhhbllnkvth6ZqYiKLBQK3TDICcdd7AMVANIQli5+
xIeoN1X9pzQxyvcczwYkmf24Ifnk5kEjNbsRLYFBECr0XkjSV5bkLBAstFnCyYKn
mJgdGeqef6Fj93/yvrD/sVQxYN975mvLLjxzCOLVKw79eeLxONZ1ifD5qYxtU2hs
mMKiKAn73em8lN9mfbPVHaRhT5wf97QAyV0Z9sjaY0fDn9rlUaGr05RJ13w+fxH1
hk1rYSigHH9Chn7Klh4ORD27qs1YgrTzK0I65EjwjwWZu/EEBn5O1bkMg3vzsWTu
yQIAsUc5WkHVjI8hDyE5LNQMe4+LLaon/M4a4u1eYHZfK3C+Q9rsHZWq42ouDYAt
e/QH/QXSIPA5Th2tx32h4bYJzVUFbyPSGrz9LWCe98IPBJCnMX+ZPbHf/qW2UG5H
J2eKSxF9LKML+PHeqk1BpspOykuB/0Kvbvl+re4PQ5CBF7RG5j0sYYpNpayps2YQ
6Tl33cUDq13zeHT55JVNOs4MnMJFPJ6bU4jcNJ2vkS7kJkH6lUQxE54qUA0oAA+K
ctkKsHu4/jcX7r1CSCWyB0y8U17kdXhLomv1PksnPk95yIIHKoidMiHxFrgR9VyW
4d6acuoPMUD+YV0y6pkmUxWQyQdE7m75MdjHNRMUWWTYWYtHb3O8pUDQJIH2P5wM
HGYQHAcuu+OsSKz8TzXg9Yu2+aYZYogG4fAFnNBizNn6Xi4cY0BWeESgv+GKey3s
uJ2iXTms4DiejIi3kvA1QI6vGtYgreyLFRsAhSmCMPy1yhoIpKavVhpqi6zkYohF
bJxmKp5zHgn56eGWap/0X4QYvvAJQq+LZiXoi/bzrG06jvrGBUL493lEI0efg0aZ
71VhQxW4u34Cc1WoJNfRxwNBnUAsThFTTNQJdsk3zMqnYRfZYxDzbEhQcKSZzvPV
+52IgpACWdCsKZXQOt2vYGSvPAubc54QrFBHhjD5UmVja09eWvnVq4p1eargFz1m
XNMtUpOQoTbxSurC+R5hgq7XLxHM5Bl1GEyYxFN4C9qKuVf52FoCumPKmxfYom42
bVFm2dgon+ic73VqrHOUbHtuCS5TLAXZRHrQTkIrHJUes6zPtAXd4AFGPbbBNOHf
mJWLP4UEtO3xVBkbAtqYrlhNjG86flVoDurObh7z3iz5aGKkKRVPmsyu+TO8m0zT
prP/CPElFnXZqKZyDliWyu8zLoaaFQNpELDmxKqrWqnYKLU/S1Pr9rFajTlHj1Ye
r/LZSX3JO8fmAddaITKNuEBeoqwnsNCWKiQ9tdO5VHdyzDPv/bx68KaRc7dZgsWN
J0LISx5ppEAvCFhFgXizSiweBJK9KAnvQshFpqSoU8sQAGMMIy9+aZQA9S+MRjR/
sAe1TSPQBDeQ1Y4hi8gyFfOqLS8EHNbuOOtjlKUD4Q3/gSLHoDOvrvfq5c75QOjr
j8cXxwQ8Nz3r8+ooMPlrVibgANzO1wu1Xl0/7Dk6ZhwxBgok2gPtPslvX+XxJqwT
yn6hNw939EPhT2aN9mgBz4OTzmFFHZ6wK7x0cA3QsLIySKvBy+Se045bkmN/HdST
W1T7nFv8GZXdF9HF4DwF4ScYOBWMBVolFEcK1mj3s0zwPoGJXC7XaqjBjs6H2MSX
mDedetaCzap6OB03sHtu/ZpMMXDK5xd92j42rMk92vZgBxpexNeyZ6Aq9Wj2E5Pb
S2TaAhqoyn+zW2Fh+mH6mOMIYiDiUXbfNzOgVGlhmVaLi394yv78Pt+waa8kuq06
rLm4rDZZDGfLt8Smi3ysUFHLMVCi+ZkYwRtCZxGY2waHka7XaE/dgsbsxVMRBbx0
Bip7uJR2nMBB6uDgp+B2gr2Cub0qkLJbO99r3/BBWCwjD9q+TTGkean5vh5mAPJq
Jo1+2H4r7+qCdvpJweZG1z+6Z/GsyU65nkusI9zY87F7lKXEkluYA635ffMdmOgb
rAtCnoAr4WyaHE40Pfc/YN0s4Lq8I3Kg1e7U65TaiL15+y8OwnnASHXml1Vpdd4b
w32XiCZ7r77/mQTzlkwMcMR0Qn86vhb0mcNk819CYt9je7wGtIa+A2Ix2mYV/ZEs
NDsZM0z+eKQXIhPpQmy9ewSxSAzddQ79/+fRriDeEvsKOIjieSOjnoN1JGxA08kO
9WJ4toHNzMtnGONnejvTHtQ7eZJt+3C/V52ppSNUfhSJwqww9ppfBnDBLECrjGHQ
URoksj/vy5Xcrjglby9DRxuCUeZmDSkrnZUrt1NphUypcRPJqQ7jQ0E/mxvfVZV9
06VBJzD7v8TJ0mzobo/MH0PCXEQpXtAOfbzqRNxe/fL2QAXtduPVuB1PyunWGuoh
mKGzCZQw1W2fAGvafz50V/MuFtKLGTGXOiiKqp/e9FJLIaSvWHImt1j8zR8ev+lb
swj6kzFXRY1A7w9MZFIouHp2IZYm7XlpoBwphP/nfOjGdf9kyQDJZeNFPzRMq6vh
IodQ/ZropCdR73fDLQs5YKcOT2mjw439HNS5+h/Wr1be75gbJnge67eoHUKg0Qig
O9TwnS85xrLwC7Oxi5av6TVJp7YbnLdGKqjjtCikTVd3ag8WX7NsrNX69rV64szc
h5mPzritxTnMeVcQgVGYx1f+GK54hdzdEZab3Jca4HNu0KBnzqrJIowbs/OkTSaK
aBq57pvEcck39tNVNZzR/YMD/3dFifXzd0TBmUBcuV34rFVzDKnOYexl30e1qtVO
QZNrnzmad9HUY7ub/iVRFb+kVgTN1y9Shni6kbCjdPKIYsIHLINGLjefzxIKCouQ
ao6xQ5Ew8FBNTenLBLZld98PmewV+zF9+hzzu8rpectc2v5Z9+FEdjM4drXHa+QY
7EqfOpaMc+VDv+9xOUoKLFJTdrx+xBOH3Juz2cfW13VtpyDoMZebLDivP94Jd9tC
wdZZ3ZgPGztFYlSpYuUJixSd1uIpKtzCYVLFC2fkR3gfmKKp4F8Z99ic8DlpkeWz
O3s3RrxCBXjNiQ5keDWBTKSrqC2btx40RcfNYJ24O8lwFXdnW4Df2kTl3QVdBtyB
dIQQK812SbPDSuDH0THM5slRldGqLIYZIBQHQ1OyGpyuNEvkWdoQzwKEZctBwEfG
G2BMt15JcCVIXNwKn2fv3t3uh7miLrlU2xv8rs+y97J4lC6Xn9QTfViDJkcMgt+T
keFqjSLpZyI6dX92lzuG6T73JRA9TsF5xjfboUhs7DYXSGlCHKtwukLdnnU5Q0v0
FAnooL1ijfru19PdOMQngQ38+rG6NdReIjyWp4wDvaGz6tw6VZcsnZMTImfEr+8N
1oCoa9VCf/ctFtu6vDdnHRkObaJPuFvgOzs05xpuPNxN+bZL3FzMg7qnvyhAkBMS
llujcCcFPvra1wwhdlguDHuqGeIm4Ec+yUA0opuov4czSjKzHRO6D17SUVUOR54T
/2jnFh5yqLsQvWojvR569SCTh7BYxkF8Pf/1kjuaJTSL1hkuOXJR3DldVNE2LK68
BL9zfIogl4vG6BoPau3bfktgo1kWO5RLLplgqVcJUcLilsom0y9Gg6YogwKsA3Pe
E2BJ7V2CcDZqn1NvGcwAxnB9UIx9KEAOoyK7snO0T/mVOnNhpyyIVw1tkM0CUc8X
TO3DO2hlKRVCxc9POzuhy7QIhNLybsFmN2IMMemzR/y65d5Qm4tCtHMBygO2xYtg
qy8drYaqAl95lAXri2WVilaVQCIsOiiCQdTUYq1NmD1otJmfo3wveCiIDe+C2lUH
/kv59n6jQRmSK8aVP4b19aKq6OQ0jsjPOvvvlNa7K0p7bRlsAFlL5UO8KTWnCdNZ
64ChXEjFDajdn582Qkv1Hkx/HmCxsWdqiwOPNX3T+39FL6vWT3jRpaAhcKUEZTZ1
H7y0bKykINEIKAF2x87NCnS3L7JOChs59GDEkv1894OaOMPOA7nLuWNBfSpTM4fl
/bz159U95lh2yBpC2oM8cD23yBrAwmZN/wUyeZAnOr9+BrAShwADJkiy/H8+s5+k
3yTr2dWy2krD+2eY6nYQyuJbosemkex0acZkKU3wgIshZHrqd8R8Tr+cj7f1XcG6
r9k1sF7jbClNkambjN/4ZwSpQHzO88UnsyZ8gvTi0mQLkqb3QVTAyKLaz1Tz/9IQ
q4rHV5PPrLr5wzwv+jMff8zP8tztWUCruG1vJP9JX1KJNb1zRqCVDUtOggsvF3bE
rT6+qjJQwXobo6DwucZNqqjWPuXnjkhxicxrjawD5mUCBiBcJDvqucBs2kNI3fg0
fqAh9RZ3HkHb4/AjMalxIb9tC8EQgbeRB34oLDYh58ya3DQfziZIMtDWnKhe1X1H
oUV4dQuYtx+mCyzOkHWu/iOt//CZIB9LTAGqCRZs0ljtKQuntY/vD1nQ4BR4qzrB
mjRFRSnUOdavuBn2+/8zSDNSuIuZFwybEss/6ArsazaLkxdmqLvC91t2oGDnmSno
2/XcAhytMZfQ4HBV1fU0MMB3FJNbabUXHMpnKdAOWOQBmF9ofCv9ODfdegCHVre6
YBrRCmcHFsMgH/G451F+076g093Oy1UiNYVWiwy+LfhnikroP+qvPWyvtSw81d6z
HJoitxrVZfJPHichfrmBf3SckJOGQeKC6bPTC2kdXxeAG49YI6CB2OcBcC+vJX67
XPZjbFj6xKSVSMfh3hKxSCPAfqNkW6KhcT8RByN/0fQ0IhHGRCDOq9hwS7R0A2nz
C/7nHPcjnk7o7xMhpBXqg/R4kOEoXOXulefg58jLT49MYgHUx10uC+MG4qdw7Dnl
sEozEFgPYDGYdNtzFEjLSRMk4Mf/yU/uuxvB+uYXvirklZWi7L6av7RQYkZUdFft
Vcz7RIgMBdcoj7KwmdGZuImzucVwazSxqbSFstuSj6E9OZpiNUk/IOyt6akpCIZn
6fFY+1TswYBZHP6m7pYTnbNnWf726+o0+faPTnBIFqQwnsxFh5Mzgsb8vNrpD6Vb
i9SlpO/8Wg4DnXTTy7qZ/I/uT11PxnpE0HC7NK+DgMGD2lDdljX6Nij2P7M9eZVU
4ReMomzcy/s+nw4ZcqhnIItU1/SQLBJvwcQS9RGUUXX/v+wNLAPnsOg+Fj5K53mH
HGOz6xfWZotB7mEtWoIBNioM5YOink7+c/8xCzVD7uA4UY0l0UEAsWMDliKpU53P
gy56g90HlsqU23M8UHwYnXdedtGLIKg5fCn6m1+09nzPh0qkeyALVSeVJMZWc1KT
MkTWEePrCLVuoTjuAINsnVBP60RdZNOvlYAIBdQxrJEIGi0PxFFx9/kmynZ8VUHQ
Sw9dimLtSFOAecurJ2v9gMrQfY1DnGAOHKxzHDI13p7de6XgUjVbQq6Nik+cyWay
/qwwsHkdctUJDypI49VeWGPBFxVebd/AOwbTaVeowccNR8KZwxlEY44HhOEEPcgm
DMbsyDfZ+uX7k/QD3ip+f9uUN6nFlcHCXOmv767DLTFq4SQFGTuMY+YgPCT5P0jX
EPzbw6d18W4dLtyQEGaPdhy8qjRhsVYuyd5p7B//uKpskLvE+M0AIgqueeuw5R/D
EefHfbK74sly+tRRdoZMxXi+2d0iDJSCxeU+Q+HTnS+sddnYvDpFNMWwzqjX1ckq
cJL+NN0WWARx9BB6bve4c/RwzczRjhsNn1CWySJaEypPP6QTzGYarR2oTCbk2qPe
ug/xCmzl/OGroG1yksc3ifwXJ93C90p8lT0MFJCrdAWTEMQe6LvbATwOVh1Sqcfm
E91UUv2bY5blgeM14aw1pvwHnxkz71sIdmQ+u0TaAcAldnjQSgCE0DJ6jBTY3iLR
73E+xMs+bYpwum//RvCGFhStUvme6T3oCRsr7pUssVrnxJVYVdWXolqtmAN/Uevj
lsq8CGPxozTuHJ3gUj0yVqKXaTuuEic1WaqFx7PMo5ZtPClUmsysbvW3tzbBVv6u
VhHmUuG0CnINBBEyPN6JKDq/VwLXYbOa5q8ikGCIgRrWkje1DRotljj+iVFFd5rK
c4+arcfOVdYp+FRqbUOCDK2I+OnMv9amTr1kbnj1Qu3+uM61fQcZcpGuYAePC5KI
VptqCuuh3hZaO6ggkWci/euq723KnJv8Ji449CGKbDQ3aWjMGSF9E5MrVAadedo9
8uZzywMz+QMRJhl1U8GWXekTXnakxgucZPOW9eyBkCfXQ6nx8hha3Iv19bNi2xkd
tlw1zRaH+Q6rs/b2CpPPZkwb8mFU1bSGaevSiTJNNuVvWB5tcJsqgn/xf+6Dh4A6
fLLG9UpMurt5ZddZDcD6DLNu/mgwwqyYw4dMmpenkoS5/Ed9jofQvx6SSEixSgOz
/m3DdWdyU1jq0IN7WpXTmq99LLHrv7H69TT+ySjLh5DDy+n28rAORrGqo5YpAnog
Jtti0kyosGIOcL048YJ2LgDqa3L7RGzlg1IQNtlChs6JRJWBzeakplqa6kqUEdsH
QN7h9/ZKw5P01C0Xm/95/5O2D2iA/Dl7jb/bHZ0c7QvkqWIq1KUt7onHR06jPUPy
AP27Rd0nq7OG1IVFliXERj8EyjWASP945TNQNo/apoY5bvw02PkEEtS9B+OsKDVW
0SzScclBmYNXeDOY84bcboFFBgtSKsJobvLOa3YGXiCIKtLVxmy7zpRNkHrm79Rq
kIyz1Mn1oXJnjQAW7iy0k+2Wn41du7g/i1zTLsolByK1nxElpuiVw0YmjjkDirig
MH9RzNXtu+Jmq2BwgfoFrxfgnbJ4g4rT/UdOrE2FB2scXmO52XgD3M4cb2dn6TGT
qzurmqoNvlxjeSfeQy4RxSN4Xu637J0WSTKnOvTi0I5Q9k1/eC5PmItd5y3qVB4S
FAkTQhE/XjXrZiVQPyKjR8Hs9NOKMwPdRf5zJDVA6KaXVa5LHtcjf9NIAMCfAeLz
U/AiVi8RxKztJCnGS5DSiEfLP55HTcKB0MxFJ2TffzMBy75OCITC3qk31opbyCMh
yLgqtZJ/SsD+52lrOryWw6DigeXSCDbUKFHOM2xB7LhMHDZPzXJgnM6xCPH3586B
2DOyiK7/hzU8+eHrA5doBPVrlNceDbOYUcLJD7caNnwg02TGR4Ju3HujAuYi6DLW
Qnj4IRuqgcAm0nHjN1UyQjCPs7/NVmHjHNujPIvUvZL4e3EqKwjs1qk9BJGEF+A8
lUb48moNQOJ64s0EoHC/JoQgzTXz7r5QcVeml+NPO0AOG5FnzSBQixPHLPkwbelx
5g9rFaMDvcaZ4RqH045482qCpeubkP7oYLAd1UPmAr9mKlCX3z/nqs8QV4kulwTr
00KoBR8S8zvDz/AbA06+Nn/Hajk8ckcaPF7BtNy8V/KtH7jjyeG3bt5IXflywbef
zTWh3n8dSKiS0Vkr02CO0A/EWSZboYQ0uwSSXifBs1zw/LSBXs8blJgJTLgleYkf
S15T5sdlgn6QPCJ9kdOQYheiPWf030SLoUAZmmbAwnnjT26ef7b/wsDS6+5/QcB1
SlpADG/m26LKGFwgyNYaNMnlyx7wDQ1nmLXp3lyNQXPVRFc0hlIeEOs8AomU9xMv
jRSZfs9v6yd8iY44k5aFN4mLkV7xgjgTkpBZ4wRhtQjoy+1UWptzxOsU53eDfkWS
N6LDVTGDmK6P4wd8rxty1+QfYv/vf2Ym4gZOOZtCXeQxIiOkeNE7M6tgXZDKLq0S
tDFrV9s7HkhT3FFCUAzQ63jBjSwjgoANv4RA42s0r1bR/cme8huADO4S68Js7dSG
czGQvSHumlf1Vam0CCMdHURQ/fFja0Wly8BduLiopZhNW7o6WkLz4c2B1n+Woc5N
PjbpbcjTzARoh/VpaUMszuv5wLJzUNzfDGVqnyndLAgj+fMdp2T+vQByRO054Odu
DYzvyZzt7l06A4RDpPTxBejAhfxReSbZIXNFUA5RHjNZKMuLyR8MBGiqzI+Sn6eR
kdtbkRrM5hA3cg0cunw3Em7YvukRe479v3CFdZvusa9P6aoEppNgrmPuTxz2q4vR
tMsB4PgZ/FmR/RCKKCoYrmZm1vgG8c0F+CQ7HrvDqNsx8iipoAg6fpBpATNVkS/e
jxu9WV4NHmlZwylbpN7tifBYaxfevMW1WwIXiAyToVlxfiaeDT7MhKelWl2WGXrC
0UNzaaaGq9grQ3zB/s9X0YB2KAAPjM3dxX+iPuZ51oPKt7IeMQNpalKLIAnQQtf0
PQb1Mp+HVlHriDllmd2DXfwrGGcJtjM9p2Lf7y8zsiautTpEaLrpxkBFW82ZHE/h
1hVKCzelbhyJiWM6BFexe91wIDe1ZdxllLjmTNPnrHXuA++sNL27YRTCFyvRZW6H
xBMo5HBlKVR7DLJJKyf1aQKjdjGBpENE9t8CsPcuAbARYb85uWZcl91S5ZzQygHy
VwCjYFZx0YB0e43f+tVQuzQpekDBV9Q/8bWpvQIFDAG1HtFSglOj6BVP19kfakQZ
iZADHYzco1RvGu/h2SJqyehT2TJN+5sqNs0cNzcrlJVyg9rec0ijOgo+W42YJDWf
O5nWP+peUKznMYpPkpBSKkVwsDwtCBCWaaQZWCyZp3F4sAoerVRHYWUIcQIkEow+
PX5X0BYnDIerOrIpVqdWXiqczuew7C3e4Moogkw/hYvUSGyi6lP1MF91bsr+YItb
hEiEXNpS29lsSo2B4yG/cz8p/X24ZTS57un0JTpf9nLZ1+7gGlKe6Yfey66so6Zi
COPNaUrmvxekIWgK4DJEIJgNX27IMZgYIY1U3Ccp5609f8SY/Ya9Yej5SsaEY52j
o50FH2AnhCco17m7bvhScNcpNrXzmpYON6Pqw39aOpRb398xPrj8x4Jc+7bO66p8
QNHXVS5IR3z5TYpBW4Ph81VzAs802yxcd/kF8IiC/sEP/e8NOvekA6J58fcDRU+K
MXtKpbwo7Gy5jgaNqe+RTqZeN3SH5Jv8hwTFfCJuTXy3EASjuCaDqxin0zzu5+Qz
1RReYa2quLrfibYF1T+R3bG+13+51a1bkm+YObWn+GCG7YYTPm7pjJoKN02dEM4E
g6CDosyZ0N3adao2g9BPk7//JhCYCaJ5XxNv1RepiV1PoGyNMcdsw0ak6fJfdDhy
U44xOBcz17ITxt5g8UQ8px0UuULAMVIT/PBVUItyhh4a7IIc5Vy+EkXqsxMe2a5m
xIB1QZNQ+/lbJvnKuzac51L5UvH8mSyykNnpGkZ1vkYP5dRE0HwKlw7tjwM1LwHK
vcYZC375qZ2whbDFBN5ID+soPZt5hPTZVCDiU4K0yJCE5lPwPI7J9fSeBXDyfjfm
G1zn0HilEtJzjHjuiQo6+02Z5YLlxjd6EES8DXJbbSq/UbKQt2uIBRH6XrccYmS2
M6qAV1Vc7m1i/Rqm1S6NxpVhxmSXvSIEMvmZ+ehGdkxEV9KBT7L9kmmWYBph7zXa
sokWZBcBI2St7ZoTk1rYhrcqoxafCziCnvQqhL+D/bAFadRKhHbf10QHOCjwejue
I3Cp11/3itzOU7EWftN0mfcjeB3iv2itT/a/8L+0fUsmhDNa8VlEdb517TL9fuRo
gz80U15n9/lqseNU+c5RC1nvcE+e16xUF8yPd0syPITK9QVhimd0joCeJ2WcmRz4
YwWWndxkd4NHtQqSLA9l68JNcfr5sLGmDDpH6FOj6n7W/qY+2OK0llps9R1/fw8k
TXApzj06aRD91edJwND6SV1vRf6Ek+o8qWWbx/EsDPJcvLP6ioAjzdsIIf06b7gE
fS+09EgbGJyMOE9g4+Ly4LVwBH4nCWhJMSsIBngcHi73jxuuhSb4yzdHguFxEAW1
S/ydSruuKc8i4UVEh3kYyHWeeCAegzoX0FG0bYWabDZkwou6H5y3Mcy7KuzjzR4q
7TVAa85M6Hdm5cD5tfKWNYNp/bHowP/LOSeeuGc4i/IuTKdVi5nTKeTlZotyoyV3
oivNicpn7uNUOGX7p4VwymvFYky8wYdoIkZUC4zSfMG4SmQKFVbTCsMRDsL4kT3I
7qLpblf4d2Yc8Stkc24458Xh5ar1ZC4fQlLJGmlb2cJcRDU5dVwt0s8teIubQZ2g
xSakPYrFkGgla40oI40Eq/gk891o/7UVmEUum3MONtKdTcvyDWruFwFmAhQt9LRA
T36euWWfiNDOzShHe06hGSNIlRCUyCtWlxT0picTe18rds1rKtPPFVdHN1vBdSo1
sUTn2KiF1BCVfavVoyFjSOaygydhrrK3z7ONONTeeZhCVnatlyG5NryHVzFb/45O
tRJ9k1S4vLEHTu5Mb8B34Da3ZsSDqk0ACIj30l93Mok9a0gfzMoFNrHI9lyhOBZh
UiGGQW6Iog2ELfgt2I9A1XJVFVcbNPOarTrO0CyHTye51MonAQFs3JD0UaJe6yxc
8rU7FSjahs64UZf47ylP0n0ellwgZ5FqG1boH8MxkeJyKQPcumaaV9srDBDmNLLa
RQ6Lgn9rTJ4qhNWFqMXf/FQvB/2A6wi8PES3LUEAhzMBOOFKTm3q+/q0A3kz/c6z
EmGhTXwWLqiP7AFL5MQbh+NPO10Nis+9wtIB/AN5148N9Kg+lMlaEXHNe4uETcxH
aeGou9kpQOj/9snTVTJubxGycGj/XKsqm7F6PuM4AP5P/Zt4xPLzDAexHPts2tHC
zTGwHBGX9H0ljbO0aF29J90fGkdhUgiedhs1UNEDdSCPFr4JilOxnH/b8C63uE7e
DqDY6hm71S2haHXIN9T5bOjXAOnygrssKzTXUjaZDLRhbB4TqJ6B1wuSyrcO+9AB
FcF9rWuEU8PWkYcGr0d3O3DDrUUX2cduURiinOGmmw5IL4Kbz3xr3ZZNlO+JP9ij
Fg9cqLHbHfmVS/FaRMvDHPqHNpl+p90iQNipdxykRn7H/cxwFfzmXocvBFZ0I7dd
mGJn7BsI96XOWltHE3b+l9ynunPqGBjxqJ9tw8xc2cPxKeSH3iS1a/bGuB0WH+ic
LFDXeO8ZcG6TKCzFTA6n7qXch3wGB6A/kop9XVbS0H/IF6QjCS1AGFAxJAxJXO9c
XgLQUa0BsrBUp1Te28/O8NdFlr/BZPWfoJONUgEJbkKMSYkO5omHM6v4Vh/EPdAf
y5gBbHUSLXJcHw83sMwsSmU0gpM2iwAHxikz3s+wGWheanHdtCFjGo8gBxCqw3YP
KmXr235lIPMgfV4rjpLvF3f0CqaTqU+tloIEgTYIpanM7vCaiBY0azF6gmGxB87t
zZRd5cD+9WcfNGMrfYqrOIev1Bu60LTdqFRUV5KSz8G5NtUtH66NBxbqB9oY7j1U
1wVG+3ySx2ZnxFgehLOjrIdJiewaN1qK09j3zOJtgraNDXHKn7qI7Ll4ZG3H/ckq
RrEMgTMJLrSRWqw+HG95L3Q+8+5Xq7UMyDIiX53zZgR7ehHEv5tto+Hl54TnxCZG
RlOKLeafk6CAJJl2Imzt2pJgRVP9KzE6B+ieI3ZoNbBcdpYCRKIAfYxhSFY1xM0L
Wka9J+JHn6Yop3zjNkl894Efp+sXliTkjCiqUHa2F965Z8q4QW4YWw8ed7jCmu+L
Cah6nKxyx43bZjSYceZ4LVuwk6QzMg3m0PiWTBHXJux/0E2g2xkA/uPMxJES6gNb
kKACNr0EIAOsBXaEKYZHwXoZz0SqFCsR3/8EBh3ddJ/i4PsDeqmB7OiFLZFthbzR
mf51w+qtFW+xxMPjNDAGfjgjXPx6P85T8LqHzctPqWcGat2uhRA4RQYIaldQYlZ4
8BULo5abAlbXXe4IxHIfqiT0mWy5wEfzLfeSUZQntT4EyGFzpVFMRx0NEEgE0MEm
yxU3y6aIXP79cgmHrzeOkjaYUbPQ4fdbsBd8WcXIhp13rdygwkCZXm+ufpNnUvz2
a/7dNyHdyLSh5ZrSHrxXyjwLzxSteWVpdOdL1AXJeZG+t3dZs4jIQ/3bscQQWIiG
cSzod2SVbvZLngIfl9pMaJfYcmmWdFKTtDNVhSQXU76oEtj9P3Nz11+n2fqHe/II
f0fRV/v659p9ASG3nQYI44XR+fvnSEsd2mRTb6lcEKwFnuzwzPK9e2+m9E1/9xHL
iUgbLnIJIIQRwFB1fQlbPxfJGpyT+//QjScHDuUj1g4wpJO9P5a/voKbif+TpZ2t
4JkXlsXbJJ9obFv+caFmAjYEtP75z9eGAtV9Q2ffaZWkZb//dQW7rvAAZ4hb3p/8
xq9ToISJPG2tAYCndAcHoKbQYd4FiCDiaGepSfugmR4easmJ6vs8DYtNpPFqyzxg
cIGk3rBNU1dv8KUNzEVBT4qCoHubbZ+r64acYvwuHYD00U2l1IUmzij44S0SDpwv
RHpju2WWc3ckedKp/axH5OaiK4n8S2E6f5zscOGoHBSVU3kp9vtGjmFVk+9QE4E7
8tT7FkGp+QqGpiCpnibMl+T0aldV1flnd4kYNRXTuoUh1zM+rcbpWa0pa1GRaPdK
ad+HMpp8xFe0uuAEQDBPQrtSIM6sUFMNw89Q6J9mhoI84hBzt3UUnHkaxLeCw16c
5HTlOW8yU7rPmrVpFYYY+nD/nGAxO7dohng6tYLoVR2/YpbIY/B6Yrs6joUYEWWy
T6jEfpWeh7q+r2MtS4UwK9eTbuve4F4PWsUOKn6s3s1AoJ92WReOnG4hADtRsi8I
Q6dMZTYReiyIwCPwA5TSyb3B6+FqeY1zrTuFiRXlpBig3uMtxJQhhSE1nGyKklFa
WRmhOHyWb3wmqnhpmrVVkF36SmeTvpblN3mYzN4LuILUQYO5Yr8db++gHGXutybu
VD2gZnuwVcN6d3MRqJ0fz/dYds2uk0ugI+buULBIjj9CHSlLurl2RlBxWladHj19
Hnu6Jace8Y3Yu2Bx3GqMhV0Kx2pMyvoA/A7fQuKj3GqtzepxJcMRl/BvnXjFacJ6
kOriWvblKajHT3oaaS+MQ2tt1jXvxd54WAy4OWO4hYNilxRtvq+nwNCvStXBvhR3
HLdPMv7n1e64//IyXS7RYHpZh+q/8xHgPOeRTzLeI+4zA7XwPNKSt8lVM30k/QGB
JM+BX6pLrNhM0bFl96M1wreRHLtNv/zD7TnEC6Uk/FO765aa2LovTW3p9W2N59QW
3kYiPT2YxiJYy1BYrUJOS24aLM7efccOoBQazecsx9lQBF4nSen/Upfc8mGrE5f7
AU2HrLdWW2Fk1nqJYo2xwg2h155aSO6Davx/wIibb/Z80qlWQ6UZ/pUniqqx/QS/
WegN4/sWXIRLg+lkSKIswud1Bz6kT26ZnnIHJDFN9/mE0yObZKTzkIgVC3XyPFMs
SgGsJwZLlPRLXpke7uidDg3HNmV9kAbaQ4iJefR6RH+I00jf4+FVTjXvQkANad7n
2LXYdzT0MlV1NsfMH+mipfP2nmgwmjNdwAJ+d9pnJmRr8NJ5fAAGXGU+XEkrbhpC
SaiAYJwKo121jyQCyZI4ctfFng/B+tswXq97r8YKH41PNST86GliU6eIHOS0ZbWC
O8iEsN/zP16uxrsX3/HNfva5f/OAkXiwnu0soeCaM+3Cd9fAqdKb5qIFue7YT1Qs
u9plmRabCMUZ9087mrqz7egKWI/EQQZzG2lrIhtdgTly+74737zpQDSoHSvDgqnv
rwffboOtpXMqVwMV7wCLbTdPxLwF09R9ZgeEZFAsL/CH0xRcP7Elv2inbFTFbSzN
fhkT40jnMBlMCqqihl7dDGVQSGdPh8I16q0yAXhoe2PaVTIHZ+JjeWSiaK/eZMDp
Sd+SzWkI/L/8/lizczUE84LUixXg+xOKHjGY0IgqjDnTtJp3d+i/FzR75rP+Chom
2cUw0J3RiICSLS103HIZCf3fNI5T9RwDWHgC95/I5cY70hkoLYVDoH0aanflFt3S
7nOcDcBaCGJ9wu+sIxNVthX8IvTdNn4+HwQHkTKjRpuY7i7sGQbKTVbEQwwTm8F+
D1J/Z2g1dL9iWJAUCjW+3/c1/YkvLEilOCDSbaXpKHzohs42m9YZwk23xDo3WQot
q2Zh7MzIQA2N1DxAd5lLzOdHxYJAHTXc/ebS9GrqmLnlk2iNxRL/NFm2Vo9y3aTR
OyjCUvKH3RRf3Km/gvMUTKZO5A1IWNFrW9DslEdk4hsmYoCPTbBRA14aoUk5s/3d
rq8TlBuwysZxLL6tG0wL1JtaBl8mNzS9ykRR6VE51wGHZ0HOBO7oDsNxPCUYhCxp
I/jvuofYRocnv7eh/BkKUbTOI3QwlT9fHWSkK+xa5EYrEDSiCkq0ky5rQ9r2EmPO
Rn6rU4BBbxam/97NE21f8tCBvRTQAyqTwmZlk6Afn63IdmpVZ+PsRhWVxOs6X1iG
TJ5dYg5CbLan9psneale1JSvBpQoS+OTWwfDgYuMvwfYbnyN8M/dgrQvaltsK5XV
u3xxfmBs7fAuk1uZZ6ivmRnbYeijuGAfUnwvQ2TK8GW39uUxU3E3jCW+2G2H3+w2
fVHQ5oh5PkMwiS8FAFk/y1fKCUmjsdjs4thAMwd7vh0YZyDhx7rcsOPDwy1zRK1m
PNGpFgwkWRnY0OGUXjfYtLFkLONXbAUnMHI/fb3mUpCThnfe4lH88EkJHfXuLEen
qCeJjt9D0towVv+vpdQyZ8IkMMTDqjCdd4CJHzDARYLfQuA1psxySJYS77hq+Aip
3GjcHtGRzmP6k1WvbtnwyO0NnmmNMipD5TarRae4BCnlhy1eYxSXfrWCKOy3QXe4
d2SPAqO6A5bRSpdFXI17FEWpEi0DsRucXC2XSRhbD/zEo1PcspMT4XEAFQATH/6V
MmR7sr/q7mX54Edz1S7YYCA0r0QEQwtNwtx8MbHQhVkd5itwnDuzKwSkycdhfUVz
qbKEO8v0aY6otlHKrufVijyVK9ZcA+r2oEX1mgMf6Q6NpUEshNmLJ266ZWYCX2kP
cg2nvEWc95n7gxG7MpRyxjm2ah/ROBvhRUxjfbUXDaTKkMOc50Oy4f1ADH98KLl6
Tk9K9zEatdomPxJDMQ3R/GORoB7VfjeNq7NwLiekzeDS65FkzxGeCiUIK2zyUs6n
3ywwLGZJZqwtPOXhCqTUbxx7838vRZ+dlnPNsLYuIDin9G/8sKRPkOlFbCus51Qw
UoyeRe+bjCDD5oWVL+qR+L9AmwHD4jtLqjdukFP5/smsRoWBrpB/dfDMnCR717bL
zUpSANDPdod1PyehIscRwzHWsoIpij4wYj/7r1Wk1eXxBaxYVFIDqLZkGpXu6LQV
4r7FHqeYsJr+Fr86VKj3i3/VYR2hBjzHu9TwzouLc7IH81Gat0+F47T803HdFUrn
EkQMdGvS9GHo5fZfLccyIakuKLNssz5jDOeDPSQEsnom/qSAjw0YAGYd1K5dpFFG
tpoB2s4gZo71Wvu6fUElMswVvzeBZnw+trMuUFICEo0G7fnC1Pl+Ky2R+yAO10xg
Zw3SRWegTTFUpbC2QotQEykZoe3vxtZLPyToOz8sGG+9aGDMP6h9Qtwoqv5EXS+a
zLcvq21529jeZPB8zkNmFiDxYt8SAXWImAipe5e9WVrgI+Pp+GLcHqtyejDbsNB9
5Fo5kAaXgQs7+NCCoiG+AIDbL9dmO1/9HlxKhfWCemXbxJ41doNI4/e/XOy+ls0d
TPDBdZbiw5AZDO72zS+J+1w/gse3liR8AfKpLywwrUXfSvYXJ/7vR8QxHIU3CHub
rIV0kr7I9XhGG1Jur+rBpflQsE2soXySDsTCNU8r8jo02eF0V/bPohp9YGkXr0KJ
9XtcArCjOqwzzWWwIbCMAsQMxZGO70NSaPwwTSdOX3Q8/TQed3LHHlqx9WW9OMZB
EErvUiuDSAfyKbDgxnhrZxlkNt/WyrxnxSdcZ4jdQkngdGTJz2KtbOaWe7vXPLqZ
YU478EXOcZyoOk0stq4kAj/zNI/Bpua1WS8dG5dEZJGyYoICOhiWrVz8U+xhTzL1
9G+aUN+UXxpHCQTWdutmtaAfpGAA9aiMQOYWwbzr1qHl0pPnyG1gSDdW0R0oG4oM
puGs5vjk/32Bk2D2PRv1FAdwbXu+9um+M1fS7aPGn1bzdt0oe4eNGPFKB2BpCo9n
pon9m02xkBBW2BMUroY7fc1kqvw2CvZgUwRbplsz2sOC1UJHgBB6hOIvuOrwhRkG
JcRYhB/fzZbVvF1AdoAy7Sit6KjNg0nzaDokOZWqN0xSmqvkT8u/6DUgQ+XEXfgP
VdroDnhUs+D1xQAxA4as8lMrq+aKHJuOEbSeekVBd1BJURMSExxfE1c8/sd+yb5x
SuCdYBZ+U1CTDOSqUyxeXaoIlijyZQtLSTMNNnqrYVTWdlOp78jY4SKfYQ6G7pNv
djd6qLEJQkkKObfj4WH4sGbQjSzJ/hNtToBcY48F8x5CoYy1aoCAmQVYIN2EYNMq
sRf8jw+HUMNwgpDnSQ5/eo65Zde8EKIpNUXpQGKXApN2o5ESlh5+SSZmMQiJllPl
wWmvpzZ6wLgf4cGSA2UPdhDuc4kIe+XJa+BFkQlGZzI8M5/l5UtSt9ataUOvd1nl
QtqSUUdKAGg5SsOPo545QJkDHrwekOHbwObT24RkLYbz7gQx48dMkymVBjViX4GZ
ubUsPxYch8LHt+cbURaJccV9ZexesDjbWHeqkKdgO0NOG1Bcn/MFn2AMe0RVYUEP
QtZW4mTNP/sLyPRApbY4SCjxljtvDGVJnvjGq4+bALcZg/pNcrjq1ZiNsAkndpmQ
o8rQXG3cGIF7zGDLLKZwuPm2BBoJjv7qy6q6sZA2i5HL9lxzubQS+ChmWDvZH6IJ
KS2yA0bihP1A0cak8qISrxeRSYNnUUbEnqMn7JDyxiHtUL30R8FTdH3Qz3pzs02l
Ftg3pNPt9s+dTv3LU5VawsMjCqmIPmoB1evUUwIdMrPz6IycaicwRzXIrNbFP/LL
J0JQaauwvvXwnGFzTcKZjQhGpag/kROWK2VqR6jB8RdCd1L+w+RBtH+WrsqbtGv9
erx+MdtgNptDrClWwmPcDvO8cYpK2fKQXEFcYnrp4mZmOdw/PooQflw6hOuSh2tj
M98DCam8MaCx8trtKBFgAVq33qNx8zsEuLxOKYegkI+RDE6E8R1yr7/Xc7r3m8kG
4rbBq91MKOY+WEREtv06T6Gp6QmuFGR280kFCHjPvjHkzzJ9HYUVDahgPvDbJIkg
93TYUvQSi+jnnlx2qfAxiK0hmidM+NXuJFhzZrcxRKryastIbvfAFOuQnpeMUFNc
/8FtXxeBbD4nof7wAXiyC9WpNLKRLuE+ZbGuZIC1NEW7H1M4+CcpRjnLaMS0f6a9
lU0egXQ1+TckT7q+QGbrI2WFUAo3FXffVSuGRYIyPWoMcPl2pRjQmc1Uz2U/1mbM
6fdZSB8toqUsnTiWu4LDY0zb+rR0ziiNbqEufpnto2v7Gl46W+s+ZGch/ltkxspA
qnrTaplhEAHhruajnJ+w8mDVUVE8T3/ecPcDB+BIHT7MaedcdRNz10M9ZwPmie9b
ZLeFmYU77j0UIfP+1jiej18ZjgxL3UJ5Mq5f3lROqgw7++exBPFC7Q2WgmERtc87
uM0R6Xw0PCzT9TCYGf7/nrghK8r2xq39tTkNQTnKnN5PWWNvcVkgFuX/bozYIrwC
p+JW8Ai/vs/1nH1S9u0E6KJL2H9brRCozUMFeBns2xoXRjE782Y+1MCdO0QwF7/2
dhHv2eaJoAj6MIHhFrNiSJyxcJUKtb7lzTjUzFOeZITCfTy80RfBXw8SdV9AsRea
jQvzEwMeWTrYNxWa+FnWHAt+k9irzdbXUN+2Mxehy0C0LRs5drjAT3fjMhNuY2/x
Pdp0CUpVnsC1/uV//0DSCVCvnzuz2C/rHXbiHIG0us3CmYh9UkSiUg7fK7ZM4SF2
wMlsD4kpM0V2j7wn5cfuc98SN/W39KpW11vZsyUXWcZfca6un1EHeOYHmFAYRd7S
Zx1mJQfCkynLqGuFhJCd/RYqanBAN0JVCaLJAjWNsUaUU+E1NgsJVKMU/4y4JYzm
HOCWorw/RiAgZtk/cjUckcpM9SY5t30m0ftMWJGmCckGfTBGb0Bmump5SDi+TAyb
MlEeXU0t7jPIXRBmSSF0c8p0C4idSaqhjcc5VfR2POtUXVS0ARwoPrtzNyQvM5Mp
tuO8dpod+I/CSeVsXuSBYlzjAN49XUR49arjI71AqQ6G884qnZcF8n1LAnsLxXSn
/XpKKKyZfQC1Ra0xWJxTZRtHoYWjAnWag/wEFYGbXyvxK6fhzzL8iP/wY0+w+ryp
OQ5/2v+pdiRiQ3id70huXgaDc66Y2qzW8KZrG6PWc14OqeKqfVcsMQcG0qN6vW7j
tSeqsYTou2yvwVPaajGy7TAif6dtZTV7SxKzlMYnxBuQvjH0XuLdRET+HkiFzaT7
zb91G0JHuZPNYEcTwKnt4uwcJnxP4XcuHXXZxgBkO/qnVE3+2enYmN9h5rALOo3q
nDH43UdXNDRbulRdRPJrB7Oav3H7O/c7nlo5regvNZn/AALvpmQ6nTjZImIMxOno
HcBkFvu095e15cjh2IPdeLZKzGk8laMgxB3obtry829s1AgUj1YoTLJn44Diq54a
ASor18YTOiB/LHfQz5MVIWZcKBSrPpUv++7qckpDaeK1h4997QYqarQ2TSNxOUWE
Sd5Sfz7Xgp2wyMRkSAkOiPGlBGn7qLPdnUqJZrcQ9GeWUw91noeuipSL4FONkDsf
IAD2v4G5Z0iwBJcKnKftDXw9UwV1EdUpW7TNTNQ9J5B6iV+8towzIQMFNArWTpI2
x/foSsh2Ah0vt1iHYE6eLd4M6bLs1lkTvwdiyk+nxyqkiGtI21tGYI2sx6fpUrOt
o1n+PRRpLCDFc84KIhcOXt+unBTTNG9Lnri5LAKQhhynFyRhhvajUyphWWEjDoMO
iAclTi0KKsl1Kp4dl1b7sY7lwPuN2BoABuG0WYALydYwb6qKWHBEfu0Lan17eai0
utuW1a9QcoPY0RTsGlgU7R4IyZCpgyUHPhwN9weA7cqCbn0eVpEf0PsNYXGEbdmc
XVeRlPnWQYMoHhHZwG5y8wjXBMentj+VGjxFvLe/Gzlkd2qNJtTzTVmQK4RULqQ7
E/aJuqKjzyDaRua5SjPaDN4l0h7aXQVchw48pcJ23rYk3p1QKKri5t0UaXkXGmNk
ZAcVcJ4ahsSbL3xQ33ODM9Vmz73p7uiznlMnk7oovle6e9EDD4tZxoMfR2P/2EVB
krgqRv8PJN79DvVghPOdNcaYxgb+qmL7FBQ860pjTf3yO95ct+OZcQN7nESWVQQC
EmzGW3GRLsz8YC/bNv/Uah0riUXXGJDiJvPksciigrLEwwssEy73Q7wIHENMSsNr
LquGrJyO+ypr1QrAdV2Bi30aTJXp2ZREdsdZ/TI4RaJDdWyYoF0o9CHBd75xAjXW
z9OSjP7AG3OUW9q4emVZHVcV+Z4MguiPczfPnncaBQC/m8WhrokuNrIcnsPTUAmE
VozI06u8EjhlgzaZWpnrAcEazljao85QCMS7Vro0hGC6LULy6Y0RibKATnTe/z7T
NWj6SJ888dI7IdvkPswB/su2SYma5SiYfeGWJ/OsdQOq5VeAb2ssCfNEgALInV1Q
XGJxYp/Up45zY9u8b2TMnAMWa3+Kw4N3d8GuU69cZEz0QpP22SRzlpXIsiUmyCyD
3s2CqWEpAJaTJRh95hvRbuJBOJKXJbFxDEdIxFSJQyKAqpHBK81iCBCnMjM0GQCX
Rzt/ejoU5uRFyAf/3434FgHGC1VpEdg9AzWfPfEGBeiKteJG0raQH7hAp+YhKhHd
+KdgZxWs8poUsWEyCXdSnJ6zPzytSZ+1NWYpwM0Z7cRUAeziWz/4X0FnHnP/MF51
c8/058qaHeEhSlKSsPp1YH/E8/Ctppdkk0zlHtwRq/eXgvW2B+iAFAWfIGD66Qo6
Xnodje9pFFFCOQAlO8OFCQVcKKTSVnJpuDOatL/a22Q001Afsq6VIpJnHEMtvQ3C
aAeXHIyWY4swIHy0wGK4pXTWxeW2NWWitwsb50IjxKxbYxTdynBVtKdSt8KK3hEf
57F0HhK0+PWd9PKA2xHsItn9VUuuiAVF+jUEB8X/7zUODrx53GHhyAbUscm/ZGUI
1sa7hwYrGgU2xe+lvOkQ6mcG/DfRSSbNnxCOdzaidmNgl7rM/HlRd+Rys1fgXbkc
LiarRlvpF+X1BdfhpJHPVTVoBoPf/g5R3CjiErt8n1dgRYC2ShnTPEd/HD7JnS1w
7T29ZofMErQw+/iwnj9xldjnigCwAkEmoDfLLNcCeBB6sX9LTx7d3EKe3XyQFmO/
zbntD3wjXxH1bfxYpkw6UlNuU55+u28l7SPAWo01lYvoWubiQFYy0Jjnz0mzdPi+
tN/wznhfEQSXOwoXe9HcuPjolsSxC2u9AH4E7pG83+BZrFXPU+b+czUT4sGcGdv6
3CSyX7h+zES6c5acpQMAVWciCC8Vf9EYe3Wei2afX7xhqmbiJFLrKzGX4XgSBpFr
SFlFz7ome6dDKLSBmZymZ2NnQ/HEuRxDC8X3ba27inislmwhhcZBy0rhtstk5tuV
7F4Yoxp9L7Q5gBaQ+ul8t5zrq3bmJ28QKosHMoucbkVIWoHqf0jDIv0Y4Ron4AT4
DFLkLHbbZAue5GoYl5DeSAdDAkdbGDS0z/SJhm9V5Ux0q+H+0IjJnIOtVjE/dbBx
flLz6jGWA8Qk+PNldV6b3SMOWJcGDMQXReZcNqWfrD/Rx9SyrPpFm945n49nIQn6
HShVjt0DsqnWx/CJkkBm7NXozf0nP0349E+vpixF+fehvVyJiV6yrNHki/aFTip0
TvOajahd0bjO+YfWhC6LIDLyR7o49PsP9exlOBhEp6eGq6XG6r3Mg+2jAlL53/zV
z9o2P/+z8mZB9FTY5Vnafx5wNC8iuTTUAtGTBXRmMQnfS0alcxGMFGMksEl1OQCB
uzjndg45ZDgiKoAVibhH+IIC9RmRcLFWFRTFjCGUjdILzROJTH2DJm7PWgXoRxfm
FFyZqGJCw4GDdwxMbPJ5CMhL4DQ63VCj2pKCf4U5k/yLBAiVTr/AjD5YCK4FAayA
jYQEjMmq7Y9/DvO+c9jLniQpVTHTICXvJ/nA0eY0lAWVlrvBXyKOCmOT3o/ztuVV
iK7An9koOndPYLQBwXFfwXzifnOSEPAg/SXTWW/aztN0TU3AHzHvbOny1OwKWyYD
ZIfMZs0i81ozlmWkC+I6+7sadoBgrpURSgN1HyeYb6T2RFV1Kpg6Hanwh5U9qLzV
bNLEXXfk3ByFKs60aT8llhgWBqbBUq42yCOjawBRazDI7q1ifgl1lsJKNkCCW95j
HBHxVudz42IgyW2c9IK1f5/YxLtgtBFAXlHabDPqet/aqCQm+1F8dG5QbpeSDKt+
sXQYQX9rWIWNJPCou+3xrDF0I3DlK8IfVHpc2e8y1zferu/1zt9r7VrGcN5twvlr
dvA8lKp+EsKQcFhBRNjCytBm7lY1Hbz1G3VkYGBwGSsjwPx76VpPcGDCMcfHMf1W
8JbfhfznduWxPTKtg0h9DqB9Z1lwWaoRS/b5/2QyYTIn/9yI1k4qnA/HlxOFrfop
i607AJlNb5zOZTnXplfM715nXTyT127hGCL8zj4XznDXM0kxlq/cW5pgeNFsp77r
p6vDeIfVd8VWg3JCho6OxAy+4bS8cJgkLuYqiM2s1rsnGbyFCqMCcw6HTgAtYpiI
Ai2tJEKBOvPoMvYU3yGIjdQCf+1pzwbymdeUnqV9atTpV6B+SBx1oEXq+5rU70lH
XwVpiDhGiS+PVg3JstEoyJM0BZaVHww69jiT5JtSwh5FdFY6mgyS4Sd6micXjbYB
miX7OuZ0LxAYH7I9CtDX9bYILke1RgTAAvs3zIfpbqjb2QRI2y5XOqDoZtTKozB4
IzQijS6GYT50oQbT1l/XHFgtsYshfKt3fnBdEcCE9zc=
`protect end_protected