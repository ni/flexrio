`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 3888 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eislOGByxcl/gRn8UziAa+H
mjgbsd36EQO5Ail/O6Xu+Sk/DKnJA3plA6MAfAy61TdNvxPHkCFqD9Hz0jDBQVx3
pmFj+nNWmgo0wYx89FQeD1yjTBpVLJJDbAui3tiBu15qmNt1H+FQhIMyBydeDEky
Azr68Qh9UpbxphRiM57nlhEEbKJUYeJoau9tTK/97kWR+YQLvas4BYqId9CZ7YF2
/txgjfX8oWt1YlFd5ofVvHjexTWmW4yqbQlScZxD3RhTDjM5hZedjV2k1kW2EB5U
yvDdBGo3M6W/7V2IvRu5uIL16fhGAni2x0M/mRphfvyn+Q/nVleog1RKH0hP1dYu
LzJwsf4hQBaeox8cRerrXVgPOK3L4pV3H9kotb5Y0D1OKXztFw4URePjzTuQHP2W
+uBGwQGrCwUzCtuyqmRa1e9Dua03BZR81ST3lB2ngSh4e4f7G3q1oUsrxJoXZHaZ
vCoz+2elj+nJGSV3RGBATQvYWFzGvxa0hXqnTInbyms2ZPNZ0fEy3zDs2bPc4rri
HIuM+9cQ4uNrN7TTIY/HrXDvWp5YdSD3c5UYOLC2ZNTsIKTaRKJrWaNjmM02UKtW
pzqBxZG5nFQYyi2RMPrEuCf5i6vA0MfAXIzv1xagIsSrn/50rJPlDcIko3kPh2zK
/V5evjtlk5CjlWOIHKlVqWSEzIKXttBUwXyNCd30+O9C/ryo34vVD/iU4PuVt6YD
74Cztl1/aATgRSW1dRgrS4lfIsr+nptwnqtd22KN5xn9uoiDNumK2LWtELiqfnEG
IEZej/CvnOYmKx32HDfsdcb8cEkJgDVPsmb+wp9dpBx/m+O+FrRgnzM4eDppRPQV
RFaEl1Rkk1TohA+p5fCHzZS5FCb9EGZv24M0AlX2oqqrR6U6fJUD00mosK80sAuT
1c6tHRaNE3+/Q5axBUIU6Q3hIx78bQmxLrT3HVsO3A2a2uKXapQ73wKphNwdpEJl
u2cIFXzeDhnIXIRsiM5Ly3YEkjpzS1dS+XRw5AqfVZ1qPDFl3pLKubKaL/KNoagw
pKWOePM1RR1onzQQwWjfiir+NqVl/7DIjt71n4TSf/iOS0Snp13uzrzzFqrTaKiu
V01JVgZIs9tA7O7HN1c011enUZOoq2fpr2RAisiyHp+sMvYA5aPPYMmlzu7TdbRR
4QgU8ZDf3PiSAih1gMWYM1ZoIXk0Iypggy3lw+ffs8ndFktYf+9nrRtOgiDKovr8
EPhDDjJTqZnT2rpgdk2Ud0j+USdxvlAFOResnPx27yOsZMZaeFPyhL49JI3p4jww
IIzHl3KO/oZWIOg3kYsr6YhaOFGzMInjhrs+Ttv8BDn0ebWvxS4oePmx4L0rhP8M
+WATjQWg7b5Rf2QSxr1wLQH0ZEChP4Is+OyL/8IWDUz3gY0K+RPUS7gvxS84JOOw
t1fhbR1xMB58vpzmxuXSq6aG7fvgYnJhcjCmRjX1fSPrMM+idhSSuNTXWwBEaocq
Ug99c+rEj8AQYzXG83WpIBFsVRimtUTA/P2oWx4e/1KAb1lygQYfQZje7PEU8YmD
18+Yc+XnE4MB7zcMbACXAGgii3WoCRFYqDipHxkg2VWk55QoTev5bBpjeSl6UZI3
F4o9PxegEKyZ2yREuvvG2Sk9ZrudgVm3vQTVvntQ6NIbqlo3ewJVuumc1L2IrIdj
lADUbelJVKTo94p6G1TLyrITa5nLjIVHbG4biTNtq96ZGZVHC3UdngK7J/aBCYyw
9dREOa7dDFmkeiM95MZV7A4vk5sNu5jKXuL3iNzXmdxtGTynSofp6l5Zu0CgbUZ0
j8ISea1LOj6wgnt6X+/N4tTSc6eywbCgnJSi58NY4q8ZbbTzqVnkD+4iPLDpuicK
w7tEO2dQHqXsboAAwN8lsRj5+/fJ9dglyPG2zsyde7liYKodPRvw+I9GdbOo/aUy
pqb6Kf6QWaV6g/BBmRambjM2YGii99Fr8jerIO5Taqh8m6XZIWOaZyYGwI6C2CFn
EcqT6JweS8aijOTg1262pTh4z1CpGDwYmRqA45Gda9nMgZtOY6jecj+wkR/icxCe
1OHiDqL+56DBrFDVa6J1+Dr5y09EAUf/d41sOp5q7y2sVN7K++zXyN9WqBLyB3vV
k9Xddi3JAx7CukwK0zbWN5whgWaXWRJC+jf3Ed/1UnLhROfxHp00+8ou/d9yifm6
duEJ92yHcEp0o/TX4u3RW85WRMDqzMN+UvR9F253KUGdSHdnGNCn0LLjdn9Vx9Kj
pLXG/SHClVr9d6i9yaFa/pJst6Yzz1BjkUNUySI7GMjrRo3vgoQEK4sulxe4y3K1
+UDIYndLXtgr0MkW03cSGWzipbSKFLzUPpA/9WyUX2j+363+SYP2uMNtCr/fHygm
Fra8GRNPnytKHfiI2PWIDEz1R1Sk8S7am1Knno8bNaJhREX9+zwrek7f5zoLp1PV
qgo4nfx1xoDmZpDnddIXRrZfR+KnNpLx7J0JvnEexshyaepEhZqIEta/Q0PWBylN
We7ApLe6nQEfxNh7wdUXd1wOF6X2Zsml9ZlIrDRWQUvxz1gLIuOfwNSxLfm4KdAo
P98m/wTJ/f+Q8keciBhGG1TGR6WiPXpwB+Cv1Ol4LWzlTPHiIGyUeEJdFB8Qg1qI
PeHZaT7ObafbIPMwOBZ+qVG3AVBsK7gLxHAlZIjBTb84NyzMjHmmNfYpUnlWtqt5
kBLuHRDXyqyex2CMD219yJMlFxvydI3rsy2eHtrYL+8lskrs9zQryWl9JssIIv84
EUMfhy8z9xYlojiF23EzzsgNuQ44F4vsndO/kApNX6AdCfr7PDGcQ+vgOQCbuznu
zKYswr3rUqGY1rKwEMBv0xXNyLF12yTnvLiVl3Q6yGL5UvLT+QqY0XHqWcfZuO8/
7QWLzM2Qa83iElc3Uf3GbHIRZBTaRqSU2hnUgrivga0BXvapFGyVp4h8EWM22VEm
TV4+IDYwfpErO0vfnKLdwPaMf1PonWbPyFktyRMhyoBq/Z/CrN1D2XgLYbXrMZ7G
4vce61IX00IkQWbnvt6gummgnifm2B8E3uuIQQYgolXS/H9HbA+G+9IHc9U9dEdp
KKu7xS5RTEhTGiJK0AMLAhaLhWk4bWe9X7UKMnS7eZAa9G69/ZbrT0chvwsT1AQW
1eKLiIYU4SMwp9iO/MAK2QyPvt4YKYdGhLBOVm0v+he5oYq2L/xkr4arHuwyHHqa
p+fUM4vkinlZvsBVx2Ja4224Hz4RnRLzmutyYyQGiL16HsDUznrjoSXMaI60vJxF
D0SabU2kLIAktpc6UDCYdndIF5kTyTTHk4J9IELbiaYtd9bZRQOLThtlgbqQ14YY
EnyjH2g90BCDbPGIJhGfSR1WcLDyHBfbD7bVtcpPmUuHtv52xO3nQt03e/B04j6Q
z8Hd2IyjkxvkPuYMDqGVM38Ug8Cvg2NexCR0pBMF4o3U6hqRcJZPOO/zJRtfruBk
yvxjCqPjSXt7IAgDYr/OUDi+k0emaLewIE7YBpeRLW4fjm3roxXIxudLTbSwMgJY
P3Kp5UfrwPa1oxgtcRGcA/YGMK4P0PKOdalAz57fkYpVF3O7V7ZqFQSDe/JMbZTI
jlDE5lPxECVDuE+fkt1c8wcZDIazGMBpJE9onB7Cm9BRC0roKZrm+OuovKEkUbtZ
UGXoDnlUTYpWbI07EfnCShVcYqXB8hq86BMWswX1YWBxZPSOD29xN2j16HYUb96g
jD2pPdGvYlqN85wh1ZJvDarrzWDDJy6XLQ5pxC4McWZcze9B4YY2LkZRhJxBPAOj
bNQLEJEy+CBWneuqEtsWZswndSPEP9zrr/gMTTiD5+49YCZdvI0+RSEHGJKGVJhb
FEEffyYi1JHT0vuQG/TS7kFQsgSEPKEGM9whHQG7VymJe8O9BVF2+ESNYZcdiDur
IV3ZAgyOXWDgC4LMYQ0c+glyApB4oaOzmxv2JuVZO274T7dYHJDuSzpv9+T6PWZ8
DXDuC0QjD4+GGIK4mC/ge94GjqUKAkovUEwBjev/qvm+wmhAUXNA4oMxhQ/LWuE4
Wf87XTf6ca7ctrlq0h0IlhDf7qupQBAkEDrdopsk4rmDc81iysLI5fC9mmOY/0TI
80dQQh/uZ4UbdvUk+das5SOeNDgCUFx4/B92Me5j5EFcJt2L0JKgdpUztGOplPMG
bTau8WaB5NoZva9LiVKTSKFIYn1z+HuKditGAgEEPW0uEm4y22pT7luW+a2uQent
ukw25Ld6zwCBR5UewA2AnkXvEBqH5ceeWQ0EogjeK2qxM01uHjcn6DGwwLSsqV+F
aJOzRrAlG7KeEzd//yxDb/UXNUyOaAfiLAvqe2fC/Bhy6m+Iehz7FngJpwi7gSl2
SvED/0gWgISelk2Ctsz2k6kwHtD29cclIzRHeOyCZhcYLSI/cJPH+o6DV+9AuS1q
26VNQTKfV//AfdP69gHN5C5gBrRurpxjOujqtCjeUyHLu5T8WrYgrg08EuZpsmB4
4y8dnonpUnRUKUeB0BMFgddCYs10N+xFPLZHJNYgr9nCKH7KPb8g8iaqTzZNlCR+
LYVxkjvZaznIWSfRKaREkeXxX1QG++Bkhk6Ux5P61v9XmEdR1+m4V1pVktmuE+Bf
w7/EBv7Jaz5rlefVlTbb43OE691aVgag2axKzaEnDjRc1AdKmshZgBF8XHWJMjDY
T+pPL+WQ3kzGPU9YDSd8UMFrRjQfxaVXZcRkCl6GmL6Hqq2Nis2BiLnglVO01wMG
mVya6VAmVU/VuhF3xSqEp6jVqmG8DSP/Q1LlVkv40UXR9JLBesWqZXI1U51dT9QX
9W+Fx8YeCLONZBhc/ER2HuNa4+UNCONyt08IzypSkM7WwRSJI3IpgLcoZdLog3Wq
Y5jlYpfhK2Kjc6Y+fveVX2PpkFPjTfwUxpNPMjKYx/ulKgPeafClkmv3/2wSVxAY
HjlNIRX7inwpkgOYc0zxZdd5/aPk+Jx0cwqpp0a64ReMpH1o/qZgOTpN9DF1O5tb
5Ty7pW6wFfjEzGDL9vIyK6KMWL1A1eHKvmhT/rBVRKSKmGI2JtsRrbfxF68xmJIe
`protect end_protected