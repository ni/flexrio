`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 1952 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
Hlvy6H2zfj4AUHTyg3DBV6SusYNG65epqAFIzTI0ZG4rqmUTseRohY0RaJZORG2h
SNefE1J9vQwpTRJq4zyBMPU+0DtV2WrK/qsUQoXCFLdXEcxdSbhQ/07fdPOw+36t
SWof143oEMpXXBfevFqYL3cuvTTaZCJ7uchQkAdjYQN/hE17s+Qjy7sEdvacLeCn
oUluNJ5s48J86JPp5CDiGQDq42TD1ZNvg89ByzcLe3PhcELj/7cjM2HDL37e5DK9
qKIkKywAhbRYZlF84EH2gVr/Jm/Doq4XqpZd7KWk687mnBolCT7gJOSyEpMvp4hz
YBo4+uNAXFi8gzOGHUTf430s1MNQO2xELrA/TC+z7XwzqZVkU5L9CdB6UxgZrBGR
tMV/EvL3FmlVbXtKGjhiI+LWy+ebrt/Nb5jfcK+VIVRJ1jn1emNe6rK3E/Cu+yB3
rRfyAJhQ5Jbk0spHXm/eVckzty28RfkO6+wpnaQ3sBOnZpPjX0DNmBM82+RCb7z5
SJLUsrvHf8vlfWPRVQMijtcZSek+I57GArciGWMBzpJqJb3qv8S2w+OThCgfrqtd
Dun6iPmnGrtCTxVIKaj0MOREKitjAkbOwi+qoXQPGjMip4hUeurF7hdNkMrWi6fE
n6kq9KX0xHlujIrYncd21CxxIiUmwIVDV7ZJpw0akIy1aRP6ZL5wlk3wvBkshwWs
L9A3Pv4W63lgCfv9AI5GzAHVnhoYwXZA6EAeFRgE/t3cNftimYoRogeFBobPnSOx
hMmgC9HAACWmJpryA+6mTgfIDytJzEamqirXreSR2izs+m0JpqUwsirGXN8MFlCz
Cj3fyyl+sqI5lu1oKN/XDgvZDI+vFCTPYXwQyV02pOYDXzqbs4vzTbVH3BEj2fJW
H8ndYWbaPZcA1sZqq9AB8R+uU7klG/x4BxMYvHwdzlaiRoiTeZ01OBfwOuHTvs47
9l2l++aNN1dKw61IdHO42eO4zCxRH7JqhZLGgfUil8OBSuLCSE+nIRUXZJZb6xH4
70PLVlLxavYqcoOzLvlwFYMulbMuurjT2en+w/1aBnTDq5bpBV/hZn9y5nRfk1r+
TY8dL8JdTnLSJ52bBJYejfMWKPY1vsAn1MSj9LHi51IcDicDGtbQS4zKYzwC8y82
HXNCyaX42kyPS4mk6/0yBWFjBz1MftbY/YSHauwdbmmy8YRdQSbvuUdxUA/Jx80n
3SE2/M1Q/TgCZgRCJlTxRCV2313ZyDRIrg0Fb6Pq6FOmlmgT6uKeKQhhIUyJ02uH
ocUIFtRJsyQy+c9Cw609HuJa9xzhrYE8CLnGfkEWgR2yVw2wwla1C69O+3ejlH3f
Q+3S5rFpRrrE0UxErbEn4Da3xFixAFN8f/a229oFCPBduToCofMZPE0V5PDxQqf1
kEcjP8nQRBuxtZ5xcaXAMrBHRw1bJNjs5SfFjr5Z1BXhmnaMwLglLAt5HQXVST+4
deqds8u8lTjO//ujKu9rrviisS4oAeOx7Xtb+WAUu8cOb2VZOeUngEXAE4osW8Gy
xerkXPeQREUC62bf5pDheUWeQEG7ssRCt0g40+QonLCJuBq4Wbp8654vBpCeXm/W
DwA2ZzLz1rqWvCZeTw+iqVDixfZuGxHkr8TPY3QKbu81J/BT7kzJ3UR5PSaL1KYt
/tQsNNClPldzQY+qaIhs6uCHfrh54Bgurr/Qh6sLW2S8SM/eVlB575W+9JtxuwBM
O71vbBVSIbaoce2bHxb8pUC4WcMZW2Q8dILDlzqhgPPexrdOS3szKWppGS9SMMbv
soLrhompD+3nQGmACYf9gThB3woMLoPUw/+SxwYiD9QUgVlUfax2pxj9UBfMak3e
N1xBzO91S5Kgw6i/4Kxs96G4r/GSfDv6YWSt1mMHCtvkiqsAGIx/vvtRrHy3N8cC
WK1ZcLTeTiePbsqp3ji3hRSAGTFEBMzAmGvhZMg4dNMZtcOH4aS8FKTcnnokcPpS
vbPj2D2wnH0NYjezr/I4/gPUK8L/MWi5rNQBOW2Y5NkwduDO/wBeOphx8xq3/dj+
ZTag6OoL/dbX0/nKyvttL2tkXNHqyLAYy/myAq+kahSB1BLPJ/ddExadH79qwHwk
jL4hIWu7b0mXaf2dmoA5wnkvcsjslWKldd+G38zGHv7OXmA1x/q9e7hTIY9/wiFZ
OkrSV8OUIPYE/5nxMD89QQsw+OC5L1Kkwq3SFGjSOUuwlEjeS0RdxaHV1vqrKIfQ
PD+3qRwVZEU3K8WQBC878I6nQmzhK76xSlVCWmqG8hIafV/wUzcR5Av65566vv8L
KIe5hxqjEdLj31/a9E0cG152T2UIAOKhw+RMx6M3CO883oGyejNGH3aECqABRHmV
oPuMcRnalkdx3VFDcHVowxK/+J659KAUWTiYkYN8vS9KvJ1SA8Eq4D1FCGuNJbJv
1cEG6uG+9PhVYinhXZ/uf8Ydr+cVEjCkH4+G8L11OmM=
`protect end_protected