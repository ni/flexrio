`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14192 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
S993bpJjwxtMDn0RNN54XzRqn8HeK8t/Cy1jDqZNdl1saeJzD7NRUnBy1GVniSZZ
bDsWKmknPNIgzn8FoPgWmpgUFgynxkqSFPGO4NueRBGOevJWhiuAxhvcW+QS5lm5
jP1zCp604FAR54UnEGVLxTCmPcTVSMqyAndbtEjYFoCW645r88oO0xORAmyCIaID
7DlOS8ojkPP/c1XpUU4bdF7gKSujlGQmCYercb3B1c3pzjUkme6mXN1QvRdkpqgY
SdzlYc8WY86CTAX/EvoLCBwYq8W/5Sz8ABzJGrQr67QYdfGr7G9+pwREweEd4cn7
OD07PhkzmO/c88Sbnr1lReFhiisXpuYli2ZiXR/fraFfCHj5A+paBl84VPN/nk59
+SMsQuE/KFO0nvuPpUfaTI/cUU43KhPJcXet9dk6iyKAuInffQSsF2NRqEr1OeYJ
YFDrtYHBJy7xXNGeTyBHkZXIA4twg6U2X22npLU3FDi3gJK5d4ngVF+9pXLoGiQD
ReeCP4OGCgjYNjac1ZBRd3AM8bqLME+wCTwZnwKNym4ozeJjs4SyZHcLbFJL3+GV
MdgMEmKYD1mnB28nbgKiXokXkgEwSrG/F/Jddu2OhCzKCDQJlekAOuj14s2W6sBm
//y3zgqpk/zSUcc63McLv+9F5MkC1EqYaKHfa4QAOo4SUvASxXHLMUsV8aL9W3h1
rY0AsLElo7Gf5tw+Vdjb+fhQHSqDDv13KK5nNhczGUWVvKUPczpjV1f+04dTiMjs
43C7MZCIPQ5dYay9PPlidjLN5WSajPIHCorPb0IlXKj6uztRyq+V2mEyCDPYLrbh
WPok2J9V7XECM6YhRDsSEcK539G6fz8pB1OzRoARZP37MlFC60h/f2TwYe3ruPY0
tygbDW48XI24eRpmfCaJHzbT457fOvdvi7tOv+gcDxiEgGu6WD/gSJicynSpKEs1
u8pKcxeBdG5kcKTxG4Rz1TpriZ4VwdLX9GozYA6rVmPkScJTsmdC0i9HgIPc4uCk
7mjOA5ceoFI/DAzxpCfQVQa5Rr3jceYn8I0HzktGYWS2McxGd9fMvoTpis5rOYJs
6EUcMGnLF88Zr65PHRcc26ccwc+Dci+a+4gs5tuSGIQUdDv/BFYU46asQnX3FbPm
oaUUkzYCFZc0PECXxs4ZfOOciGun4QV5IbgWX4cXEvX83dB4l+MDiNhwyCausgaF
P867HaGUYH2ZFbIYuBVAkcQ0WhxaQ8nM/be/7L21lt3mRmdwXcYps+T61RJb9pRT
PeOyyQU+cYWU+XixGDLPBiIKkaaKAhB1oJw5hmZWYh8tYe5yoS9T05kFxGwruhDR
dWAqAKQabO0ze/2sE3OfIWvU1vjPPD9MX/CKnvvTXSrMg4U6aywj4z3N5sanjd2t
DJr/O1+fDFB5WxmYElSiwI5toZxK5Y7ip4U1exuThEGy1bUPPTtyN++54FMhMKAD
WIHIvRTk2Ig/LQ7BGvQb6SS2mut5PwXQTNOeKOyreuLwcO3P9MCAYysUCZUxwJ8V
cZmh0uvNFh7GzgGZLn/LFAIeSZgyZjmNQp5jcgxNDd5eTzN6HKEaXA95FF3ZFWts
RAPcHEXUxgj/zVY7QykL4dzZdxJq1SE9/S4VgnUyheFNQ3wZ4MhhJUXQSfpFsMXo
SYwk5UAL1LhtL04wQRgVr5Zgsl6MdyTrwa12LVhO98zMbfJK/vv4Dp8pBEJrlIwo
3MUdD0ezlaqHxhrZ+FhW3EQwH/YMBt2x0oOE1lJvX+7XNWm/IPnruRqksI5WyNZ6
HGtCsap6w47g67OK7lqxS60efhuLXDPoy2sbHCXNOor0XMjTCUT1Ivul7jPcWj/o
jchBesgFh5m+Ql7vfIqW4wQUqa+QWI98G3KozRXAnnDvWibWCPlQl4+4dqCplCVg
B2D9q1XRhuB9ejdiEYh76bMmd9nOjuvk26YH+BV8rxeYNlwHcEvlkwoEj9yzbhpT
ATb7AxAL2lrQvTq2vH7wpwvXdSFK1xw2rRWrbxJV9nMYojNrV3/1c6DVU5TMHsXw
05tLQfILwOq/j6Uu8Z89SwFOsXg0DWH5xBNjboB13ZeJvfAhTbQHafxpbwbhvgAW
Eq6moWvE9yni3QiqQVkw1olFvP4qFaWgrzpWCpQzgKoC4gki5b4WKKVukKhEJai0
ef+ewU622RiUWZwIpYs0rVxVwEjANvWvOZHA6VqwOuN1HXl32bpy2O7jv4gnewzY
ZIaPOnnW36aa9xsY5jbHA+xiCTAS1+cQP+QrDFdMwhBDWK5y/H7QLIiXHoWImJGd
Z3c6X87AbMGZ+WI3bRuf0LjvCoyV9ikp/wd/RyOl5bkNYf3zw3mTR0MauytTcwhB
19RJ+BkuDEhQ73pGynEoXQ3IE5LZXMM2cT0BpZLHQixjWllkBB0diNOBBjqlt0x9
59HQMxGXZG0+IpMwV/38915f15sd+16vpU3HqHpDEszo7SsI2c/qEYk27OpJYw1M
WRmzzUjIGg39TETDnegqZtSmSt4R9HlxpnW1LCATY24rFwmwe9y/uzK9sSl4z3go
o2KJWJL8w5eLm16FOPDCectfsM2vujsAsXFZ7Rva8F/X2rXgvEca/SGmxT3sTVbk
R4Hxwt4c4yb0579HypWSj6oBliJBMwpr60GIshkDw3BiJ7fqKxG1Gqj9MLUk+Xsl
Y+W6j075EOCgnWKed494sIRB6rz0h9HDAkGjxCZb7Kll6Hvvk28ufhqqmCj3Px0W
NwKHhPuRlYVjTszMX4yKE1FiPM16+5VE4RkZKED2s0oSgmARkCJGTJmquHbm40vW
oqOA6UUJgqTu6bEUJ6EtY27LAq1PQ22GYQNrLX68211e3CGXjQFsCG3OezTlzPs4
TuY2Aewdr3k48jY4xH8kE18ncxamL0KaHzZVirW8dSW7SUhZpvAzFc/s21ue2n2J
e1tsZfWAGKY2Lk+hD7lzo4Q/nY3a+741eZTRKwusXxql9OGTyD0OWy6fYl/EDy3i
pvL+c8yTibL81v4uI7AkhI0pzPfsn9ArrCY4LFASaWQCfHJfMwJgr9/Qz/Yz6izt
PavpquO35ya5nXqLSZkd+rfXZ9r7hYv9uEsfYnwQfBYw960lnp7cxqmxdk2Lyys1
Ort9yiFPkbrcajfg8G/0gxEFEGiqla4xbyrCD+OujXFwbsJYdY6WqTg6OXlcPhqa
awrvmW2aN20opdX3M+X+GssnKpIjfAKcqcOecMcOpjxMGL1OOrgxSVrZLA12a5M4
rCbzzRyoD7tsnmgesz4b1Hoa2j82sz6Tim75s7fswvPVNsHOdpqAs8AfiYrTywkZ
Jv+mojWydZ0NpC8QHLPEXrsAQp/+/vQiGxeP3orVAMYCAXNdlO19TEiiFNij9Edw
7wa4k43W07wI7UjBEq+B/EWHUAybCKliEkOSeFMN/6AHOiXXrC7lXL+gngQ52kVu
VUrVNO3b/Do8SIJCs2NCzF4WwaTVSNisGlrF/BLlf4wVPhj1KxLsGaqfY/OFKxM2
T4Bk6GVNblVAXEF7qx6ZoMjCBvtZbIVzb3AKiq3zBwLq1YdiGCUpieV3SSx+due7
9w0q/5LQHgKyzASzu0zQnG0YZ/z7mZMAoVXIdy67aIVndJf1lGoB1qmLAvaukvdm
QzztvrH1ARqlHCnr9Hj3I1EoMwOe+830vBIdaxGgfi/0plsjxSf4FG84JHcS19hZ
sBNlj1Of3LuxNdF904XSnG2k9A0MxzpFxFSNuZBcW7GavNfGz7fkbJ5KuHCzU9HM
ueN1wewV/4p3sbCc6bOD/JLGdvuc0POGKGV+EuZBFaGnURZc+hUpVFk4heDE0ROY
+UgrfstwORRjtCCgxWKN+pI4WzssYFeIFlxYzm5D/lHq5dnwttU6/BpEZ+R78PUU
pFRJXLvRtdo85sPmwQgWFc3iS77afx+yigQAWd6uW4wmeMMiA2SpK+1dhNG559++
b2ZKkKRuG5+ZclTuTvaZct1oAw5xyxHJPHfakjl4mHK72FflaI0hhBrqEqw6Yy4O
txbTxFVx+r0r4zh8x28/W5PsG549kEvIsm4xax33b0CUq1fkOc7XVnsAA07mLLiP
HU63zoubAFeGej02cnCc2kDu4t5DVThf2brpHLd02XrdzLdRiNwlyW1RhjL5bUbd
eMFbfSdzRAQgISxgCD2diCRJeSadzAV0gwTC3Gsr2dm3cCXKasV9S9HktrJHASDC
BkXQtvcrxVujCaXDnDFdUmeSFPFXG+cNkr8NhyfzI2bUGVuYxfvorvBBRQMTSbB9
zv5J+Z/XdPn+MHNFX4+sDRpIjYNWAOXsso0FlaRtBfc1w0rhrObkwpCeUCrv25eR
pizTuHYu3JF76hB4c9abKlmyZYR5YZ0ARwhMWPVhlDdu5KpCrgfMdZjamxPizPxw
mhBb09rQOCL+3CTASY1/RivD3RELS0LDUK/zgVb41Y6YlkAF7NGaOmhY3WoPnLIJ
18mTcPSlxxxsFNAs3Jry1Lbdls3SxUx9+5ns9XZutjUdDFcsbIVUaNJNZxiaCtZs
bmVGpEmsHTdxeXZb3hdujzJmMB44j9rKotycqKNr6Zb5JN8RwSOR9cCiyx871UKZ
r9Wt17eSl4sWQNLU54T3CPTMoTEYjyBpAhS0XMuVO5b0x3i1v4Fjq3RR1PaIriPg
j7JDBLY+3Ewy5eQjeHplqHWHljByrYWl8yvN45q+4STK8j90VHOKochw0WsDzp5m
eGL0Z3Ij+C+Lli+fVMhmyCh+00roCQbQmcnbJPfb3pP8SymBz3Suv7Y3w4+p8CJE
4dRp2ncTWM7civm0mKbjcd/wpf6emvPdSYHK4BpVA8kxyRztZY/EL73QGGKqXjaw
deifvx9k66+lZxZP96LYptYAz5+/Cjx95Webs3iYcfEK2bvcmZC2GkNOHorAlUdt
DExpogeKa4UVIxQeNpM+ddLpCeUWJgF+JzsHcg9o+tLtcY98M8kOMdJLHJROvfvW
stwm79LOzETPVhzvIt4ojjhlSOZ++G/pNF9amH+aXhKwySUCSt/boUGonTQEn7Ku
WenVbvU5mJc1AxsCJNJJNh73BJ2dstWutoe8FnE6f/9GZn23XnKMljZ8UlyVNz6Y
X8RffFj3a+QkovgvbN9Of6wPnRtGhthvxjsMKUnurVVT2oegCzexlhhJ8CGpBU2v
uLg5VlzUYq7xp0jfS8DCGI/5+R0uHu/IQPUIMykTYTDZnbGuk/ygSBdyDbe+LSZG
WURITDqISjzhLihHM6YX4fezwi6pPWfYraJg2zLV2OlLyXlz3HZamMWfMK8Eds+L
XQPzevf/B5tRzCu9QP4XD9hB3rT/bLPxT7FnCSCD6LuPSa3QzGGgZ+9ub1MYJukt
1GmOQ2yPr+MsJlnu1pRixGEhGNaJkC0TecFYLWLWu1/eaFiKmqHoi0QQhsQiJCFB
SRmdIlnPyjkScADHgwxSue3kJfEbm1MRmMO4f2mPbamrn/BdUEBWH/oljieId7Oh
TpemRD/fG/bBH56ACgdR3yeXrcbs2s0yxUYNjcpRzK/W5B7Y7n9zFcQtz8p9vzIR
ZvIXInRSmtEiiFKb70NpGxqsw/uvmJaZ+8yCQUAYTlNQ3yIps/7ZPEN3dkPwP8ZE
3RSoslLXcp2Ak+Iw006ali5d8lowkNVudRjfKVaJDVlt+eFJJuEMQL4Hpf1zbvCc
d1LdSyn13DGYGhMK2gmlqVhRW06/jBDorSiDg6WFSYc8me5rVpZsJTDuVnIvjuhD
xe1vqxVuC0mM3q9LZ46AkFbLf4ZqBeRrS9fy+2oia9MIZuC5ZmCCw96Io4a3IfGC
AQctbM4jkOgMXFrkvKp8JyrDA4JT6YClPXFs1/6wBc3NAr1BJh1cTU6JYBQzSLiH
ri63OwWxuvT7aa3qasjaobw+2WGRBAgJoi6DKmL5Y2w24LtWJzwXDWDM5DrdwvFz
HS5AasD1vdMvDLJfFu3pbbRzgci8em9BVW3JhzpTXOwIty6Ymkm777oZ7oPJTucu
C1lJQ0OTfvN5L8NJJ8DJ0qRyUxot8/DNSlfKLfKjdoKxOXqKmbDwhRPK94uAan92
7i4gpr8T9My/lYMfGsFPoU4lqrTG5JIZS+in+tamxsKRHraXfLPuznpzz3o+WCwf
AbHFUOCP2L2vo7RHmNcrp8CuVvEVRmiJ22E/ro0CuNBU4mrFOdZQ2WNOoaL0LSyQ
P9mX1UcR7GBXu2fGKSP2dsanKMBCsMmQVanX9gD6IXetb8tNKVTJv5L8i8afDrOR
tvG1TnGauHZJ9AN9DDAJYKIIfLeV+qK5x+QjYl2V/oMdVZQTyHBBBzWipAnh8PlJ
LdyVNjpSpUJpyrp2cAplzqdX2Nqvfqj2F6y+opISHhM14mcTVatkZeG21C+cNCLF
pBbk7qajWIrmlUP5gCoH2QDqUgq7f+HdyL7XgO8ookUBMtBMJUrx2BKFQ6P6bfB2
2ABcOC1Lub7dAiaaSTDuARXvaAW6O/HokBvWYsCXW+88O5kx0fqj0uAChHf4BtoC
885YDWI/hzKnniHzSAL3DZLAqMRhjtNvKTPk7MFFSSHfbiF7DJxDLCaM8vznv8OF
afzfwAikWSN3Vuu+6WVgonx5e2SUVs6as4e6eVSiEphn322Gd5okGrq8CKtyqL4w
jG2S6wp+JLvds8nW5bMKrzTEweSIcrHeUHLYayw3th+k9MqIrfzhnRZq7mXx4Bbw
6XigMb5JRC8dP5YEEPBptHpEHiHZ4lbGFPgiHPeiEgleR1JpSAiNa35A4tdrk6It
Jt2s6BlaUxPdOYF6gD+sFMusvfrvesyhREH1sIZDiGW5+XqqCTbTpV91S45a0lgR
3LmXUIQ1RRxYnatQ1QZ4u+fwVVDh4Aapw0WkQrfL81Qh4QwP4cajom++OAHBbKiC
AGyPB7f3gC0uigGZmShwqxX2qHxThy4jT1LtkPZamy+wrgmfb3oFYZmJicskhGv4
mGlVLkueP0ONjX3hPqccMc+OvoWucyqM/AD8+DyYE35XQQV85ca7Oonc3c91bCgm
sNwoA7pGVZBXi5ZeV4s3kJycmB9oUVtXzI4NgA5JnBNfSNv/uz/GBuWWTYU2E8DQ
hdijX9onO0rzRRhNWeLczvKlO6mUJUqtlvNOvBJWA8lt63qsWHxAwbLA1fOhHq/C
gVA1XmC0oOL8UJsXtiwd6iOA894Vw8z2g336oFpAidYwjd2A78GI2z3vwM0KNVyt
WLt7NR42rCdokhTtYFN9lXCjU8DfEPxkXxgOJhymrvhKzfss22BjdW2nPFwwSug+
CDEXXUT1zj/WI2Gvui13n50F+Ol+XTfC/IES3PUizlbzRQRnUs11HFg+JWRcXUfy
7jICtdKw4Ps9lM6235dqKZa3O6QzOsjZSzQS90vRxjphBQTYZ1vQLBBO7XXTx5v8
h17wWt6YmJlmP3zUS/Z76wcMe+pB3uTZGCtpGIKYC43dNk+eQkx1p9SAEiPKNqN+
Tk2GNTv9/RYfDXSHQi5xYi7MOI2t5SX3UJsXF1YI5Yr+SZvufPfYd1J8jODVemSb
XDsCyk4pPg7BYnrtJVx5f/FW/wzWFSNhRuWKeL8Pdq9METrkealCcofwj763Ug1q
OTz/C5S0MeSF35e4xp8MT3O3jvjKmvfAQeTzVBpt3gsV9njJQfCpg9+OXK0HfGd+
otihnaLXssuUuBoCrgTxdd7eFLGIstfngwK3DJoqPqEsUBfW+VsjUuzm8ls7da+G
JMAX+EYptsKCBMnz38qWM7gYMvFdLJ+GJMqn8EtlN0me0tBuQ9d48yw7LRX8+hUa
GUCMAsuuU/3+vglRI9MGMaj6QbIKsSA1mIO5uriGjz4Nq4loGLE5iyoUv7CZj2Gn
6aYucAdnCRXkjBmYXpEhtvK7lt43NemBkJSszoVr19H7d5VsOOS+4J/g0lUfDE6k
Q/5CFK4N++puvz1jshSKbWcplrVWGjUeV1am1EwTScr5rwBRNAeIu5TJXsMeZeOJ
K241SpIc1gnOI2EAbPJ1q+xP8GRTucKsX3PUE96D5WivKFo2pYKKlTmejybWPscM
8Psrnl0quYdG97e//QryXpU+KyUUh2R53zQg/TLqq2Qfox+qAYYFWxqrcSgGQAsC
2RDY+RWcR2qLWEUyyrWET9wDM/niwuU4Gqh/H1dZTUc7YLzWgkxJxI25WPhqMYrh
a4Bb85N3fIjgh1qB4eNbQWDuojn0FU4VoNWnmYlglx9vKRrJJlB7b+uG7f8VEizm
bjesC+jqfKjY19ZNaOJNpkg3Qpo9MG4UHdcScMPZpPIH1IMeCpaK7gg/eM8FR8ea
wJ78S4yA+YNSGAUakhh2k5Liz1NCjM1CM352SNvpukEdeH/Ealbrar8Aoe6TvQZO
1+Thu4rLIfBREg2pul3u8sfRw3ONb4V6rqNLM/4kobR/Z+Lsx6ajbEGEXXeM/mcA
d4FYKbmyMfOjYo1wuGhVDWoLKWUe59YU/MEcJs8c/+nWebbOifC+5mmhhvtoWia9
rGvsnOaN1xoo8FOoy5bKXjXu4Jd7jmcEhaE70s8TiUSRvoQSvB5yh8Tw9wKb3mT3
oVPL3r+tq3VDtW4DavLEJqz6QZugJwQyWDPdFyljMOjtVSAF1hwsAaGgFI7C3Evs
CPQlsBc67ypxkPwMxDzJElNpDdpxLSuJtFtwshKxJddGYWF5va3ocbIVsjTXgcDw
xEa402Ub+mDD0tNmQaz95StWMQ+W+Ex3XP1lN9G3WlCR32MFaD+aLvylkU9OKBsF
jc7KR3o6lAtWbdxPaKQmfSdXKquxqzBbPUOfZW5KquW7CjcmjLplzsgQsQqagNt3
ppyFAl+GAR/0uMjwXOIiqav85g6Q8UhoZcp0R/qL2k2ziK+jJ42GIhgsBW0wDjMb
Ss0MyOmkpNWXZ3j/q37JmO5bsmZ/204K/SqDYWASFqYJtrKVqwaM70drTYWtHnn4
GQqYfHJHowVYhzDfFfsTdd9HW7x0bFFEfXia+JMr6B5DrA0e1eTVDUMKElO7zBi6
kmfgm2jd18r8Q2mrNbfd3xiYRANFWpZbpud/pb0HsPzKwQ7yAxO8buegq6O0V4I8
eCzEy0puE5132AvjjIf4ny1PqHsfBfTzGe+YVKkr3nfUAVBUtjcRI/bDZlcRHXDL
7RYKoGtQSMYQ0hybiMuNybGO+JEZDD/61t44gwJYkVylCITyS57mp4XbsntiSUev
3iyxSdcbcudxhVyev1s/fgk4SEt32Ebe4HGiquAB5J/6vFMF5Hu7kQhAMOp3r8sF
gQsDAli+6i4qi10w1PgGsnYvDIwkThf8rg4EB+c0UR/ae1m7M12/4bGkrtHwPaGy
tYngSuPkXyeJ1LPbkj5IdVxUDTkN1i5WnGQOA1TC7McWKFF3VxFInvEkA8rrr97o
RiW7WiQZJsFlz5qyiIfLG9uHtVTOpRIHfLeXj+kPFz7YA3Txfvd/q4TTazDMRS5U
HkjVTYX39zbv3zyLpz/2++DnJ52mxFRepp1pfDM68BLeqJid52ZSStrRVD/S51Gn
JxMpAWJ5wVhrUcyS43/7FrVYJ31Pskyw07sIbgDDfYSmfbxI70E1+JMvHZxCMet1
ZAK/ySrRPUJX+QQ0owNqqmiRFfzzUqM5zB+SXny6/4yOPcv9ySBDdBZC5QbNE0hA
OPAcVwZBZpMlAevF/6Jaa8rTbzHEHfE9dvNaTtPm9X9tYPDAA+hR/1OQymveQK5i
rUbciy+HylPLAn5i79dHliavKSxf5K8m2Y6aniBqrOh3YDiW0urezITNUlhlXub/
32JTn32rfApR4aX2D97t2kEn8f5szzQkCxfp8pyP5R8joOmUPxV2wBl/X0gE8F43
D9ZrOCBtIwRJs/o5QugpIEhmm6NAzJw1fbEvSHvZVcQDAXoK2txVqhinHwRoCc6C
PsAB6IpePw5ZU35cyvDt9Sgm/8klnSUZMh5W5PLJf25OIk9OPwFRHyG9vIr0ihQe
RwmYc3qTmTdVpONriigiQ2Q5TPL0px/PnaK7Xr69Zhc/ajfN5QXQNJcmdmD/AedW
IMCmYskFL9NDVsL64GJS6VcT1JAPrTanAKcunmfpfl7vfb+PKQdTJYrfn8A0kwXN
/czZNIklF9FkU5bJqlrJ0RVXH09BgM771no8aag9uiuCNgG2x459NhQWN4uBoV72
u610YmWqCvgaXLfOI++8J5AEBwUq891gMTC27OTis6osEk96Xd+O5AUe+G2sfTOW
ueJFuV6F+EzuJNpGssNVjHSdBKIOGvXsjumbHN8keoN1s65B7whmOO16fJOG7Np2
KJQteyg70vxhnEo5qI0TeYXfdSCnKqXiNfZ7o85XfeOnZwic3re5/L63DB+CMVeR
7Kag0L+zPmWoOsWfL2rZY3rJW1RpLFvoA18jH7uHPJM4pQJlLf6e5Tsp5GWzIVE8
iOoM7ecCWYKBmK1vU5hopdViC1PiKa07Ts9PYgKe2dfREry1imzR0N/EMbfODvtL
v6hiMfR83jNfJKQJXyRt9ps6LqJX7h5sJ0Nwspg7bkUCHeY3Y1Ytd7J2+BDOHinO
ARk+TBHP3mcH73VYau44bOOeTjR7D3yPkvTYAJYX1ER74erRHpPZEFsHtp7mLcAx
Sl3TTs3bRHaStD4FOvDiv7pgLEqt/vRxfu7D5pbEXGTDdh9BimAVATgGWrv0YVf2
XXpAn9atyXXVlpdn/uwk7/zm9WN6dNhlL2Sha6FbbbrIVpMouLhCw8J96fPuUjda
bSl4B+Gj9lYg7Kma4qw3p1tXjlb6qLolnBwOw8LOH6x42zg1VCn8e8sMWSgKr1SC
KkFz3KMpXPPMjRIs8indpzIew3xMG9IZsz/3dmDRhpMkjtJiTa67a8bCkS6AQFFM
E04Xne7GkYjU8cluOVjlFDEsgKKX8VE09ht75gQLLvCzx10g9VUImVLQ2GgNl5//
WqEDAwIx06LeNzgUW22fWfVrTNAhjo4nJF2fuC+PMtdRxtwYMyej9k98fnWkTi6G
eEGr1xafYDAbSVX+u45HMbDrqeqtpfmNA3Ov0bj2Wk1mpxqLL2DCewkZ8/QlMOXC
rGKOh4JeZM5vSpEbB4qXouIy+5g1BxOIAp9Wj91XeOO6XEaBZnEtqUDi1r01SorZ
Q0HGQFS3bGTOiax6T2KmUXiTVcYUeSpfTIqY87ufUDO6PprRtYz1jjw72+NELf92
jt3xTmCtxda7I95cyyRX/men24S2AxjDM7aKrSNzbroWOQLiAeqbjMGVrbsNAszR
b5HblgnceFcit+SaXa6cQqBMkHbspttP2jd3NHIBiFs0z4V3twzlNaEMcU42XzIV
nSB5qDCTwOz+f12XrCkFp6OklAYpjcO4t8zZtViKO/By8SM3mVpfqPjM1cvKouuH
TDO3lxCV5HN9OmFNlojhKBstGJL5FRhM47UpRnmYRr3TkMWFlN9ZkIn8gsWzrmrD
iRv/lfyfYklOW11Xo8NVQk5keL7yjk8Zq52mbrazVu/Mw8gmRHGlhg6zZe09E0CD
HEq9HCk3CTT4mRyvMQVnrxOcLK3XwXJ0gEbeSTPrP1BtFlLH2ZepqR7KCo139VZ3
+eXQ7wTltizxMfksCUXB4LobyTugmJeu9RM2zfONXA/Yu4k9zC3+uaF9bFcAOYX7
nQSenHM7xtxK06MO+leytMPl+QyaB4duiZ16koDDk9IKL8cn5xdm8w6xV2DT+7t3
wJQeVfLH8aGrkcvHLmuYbtOUTDUtf6d+0YowP8JXscs4DVw1AzN7O2a+owAFN0Sz
jlRPQvWFwqg9dhU5COFQSA0SSWrEsZmdaM1dJV+1Wo0t2KEJE2jYbn/BZljmW2PL
CA+Ag/k86GXp2OTzB2NGuHN5Fb+sn+KmuFdET3wEVVg4JiCk81cLM837ogRmEVTN
g/oNNSZHiYDatLtuW2sbr7SQvTZuCwNDQT+uwARXOPOfba8kBSsFlJxv68iqSwuf
qpUlryQT86UGdQqzZ0wGNT/ZqNqIBYi7GZgatES63C+UWXT9SDomJerVXeZrhg40
2XB73CFSy9CTMfJgoFkomzbmSZUJYdbv+8Qyx14vG0rdE+xJiFAcaC1rgjUv0Dvi
svrtKuKXwyFXWNGX4CnIShVUAdwKe1VnHUTdFvCmtAxXQ15IVcSRJ5ZRRDdsBg6G
R83JwwuWp8NQV8HttSM41XJdJedKk0OaFW/pTR2MrILr32vPfcB6Al33YqzMGMy/
zp+pFZrfF8U/bX2SjxWp2iD+UCP88/vxX1yDEWu+eviJqWJ9JLFDkTW+IA2RjBZ7
msTpCsWiGX/7wyw6bwpQkh5SJoHsmCMcQQbGG4z2Wlni6mp+IxDKKdRALcVWs8NN
AYHeP07KbWjjPXLyFTuk2MuV0YddOl6vgyNevyfxCCdz52OWx4hwZfgptfIuUSVe
ZpcaiUlo9g2JQpYuXICRQNwRqX2O2O6iZaEWnWQ9LJG8cGmg67fCfFzkL0IOx+eX
3HzlurK8hEVLwadCS676M0RRmsvuwgitDOMDH8Xoz5xuDt5RzIASFlNNVwyOkSr7
xt/hWxfdovYw0tTabECCW55UqGlnymD8FOJRvldIrMcbkwl+vLJTLyorSETxMfs3
hjTml4BI+rL/Or6x9we/osChjxuR+3Cugix81sD+EdzkIhAJJykMshVxCqwPEXxg
Bmyc2uU7rU8k4wUTkDnyvkFQWkE4NCka1cyUEkzy/eXEK14X3AYSPd+Kxh0dJ7jp
8EMmPfV0fsn2KL5MVobZGc9KiUD5Md7v3LQLFP6p5BNihfWqzcV0k5J3xqPcKtbP
hdOCjnFXqYokVt7HM8uAv3bijLkgI6kdiwQwzsYGrgKjbh2o7arLb3PtaUxcehzk
LND9BGaKwyuaBRxcLccDYUA2j4U++bgaRnbmEuGEMAgn8R7UA7ANsFRNQwMc/kCe
02A2Jdv513Z0TJ8hIJmTA7YxE5pG2BAcxwmoKZZKpmooojzx2zEy4L9cWNMf7eZL
qwRlsOhEN8jqqN77oVAuRCtOsSY0veDcwJoB4idh9IOKdmetgOtldIt+IpqYDvqf
fuddIbruQ6mscucMqpBuMpSxy1xb0Jfx/SLATrTk+jKNRoulEZdQBIlOYs2nj+Ec
TOjg7w2LBj8mNyuW0mPBh0ZM0XLEnwy0OcGqwlC0Mgh7aWE6U+8XL0b18s2KT9W8
tbwN/kOnu9yw5JJfcRGjwJNqc73H/45ELjfllDNd3oBWTNSbs/FbIMauOHpwe1CY
WoaHAFgPuh3XHExXgFCrF0cru5vzCFiQ8fRzxPyYFxI5XaYK1iepx+t+5I2PXvFL
uLFMxZHCc8WoJvAONYlQi/Mwg8z2bEzKgJ2ihhVeUN0YLzX6SeUSU4f2kSHsy7Oo
A/4wdFv9SXBq9uyYoQTmClvasvDn7Fw0SR71egp79qZ0zHLLGq0Yk9HS5O+jprHn
Wtxm572UVGSI6kA9gfORhAk+BkDgITo2htpOTdR0lNs38Ohs233QmXKYcuRD1ZfD
1GuHKstZtScmW95sviGwXY2d43PcDMnqe/RpHRtqFKKAi5qKZISM/SfRseBxcmR2
MQV03q7HUhfyKUMZNf2J0Mc+3YFDsNubf+/hmV1zdyLqRAlxGWdIvMhypt48UAUA
DxyiXFk1nLQlb7WRqGyqG1YUjajVSuMm2SrCoUird+agYXQcRtIX0wY0aqYMwUeg
Cu6hWTWk3QOaPI/bIF5o8VXUV09sFa0dGHRjfZTwD9xg1CLkKiakjrCS6t3VjvGc
TO7mHcLz8jhyzlHG4IQFsXDxlGnO2hTkV+XZJnztZjDYGLkYHWq6isvqfqKpdmwY
Bi8xztMImgXlZ3i7ueyrE52O4IGIxuQB65nhhP9aboJpCKAG5hK8z5Uq8vfsINCP
r31KE7A9nL4PgfgiCI/Y/r5F4d15QRue5Czq0m8HMZtIZ/cJjkZW7Iiz87eSj+yj
JAelssC40YtEYIVtC4EJ8C6i50u4XfkMhoIYYRU8R09PrcU7WYdDwURA06vB5oQX
CsE1jO3SsqM9O4tlLVflArEly2AlfEyHg9pCVHUZQPW0rlpBqVd7tk7qEj2BBQoy
3ksNx2b/3Wykl67bJz/FKt1A3Jvg2OX65VDhtjKTNyie8hPrkThd9dzbdCH9SvgP
wa/BlWdopEXkFhTeJt413IS/4UbpuPo0cHys9TE51RV1EbqrPVHih6JJrEYGEYEi
xX1RBruRyKjU80zCpSPEiFxM2F2UlJXKNLoNRw+OLeChvnHtRXcl3cQXoKRU2Sc7
wLu9ZbeM+Kzfv0fkHR/pmIzTrtChSeMLvr1RPwu9o9O+tRVasEZOGbDaR6nJ0Kst
E81yrOjbFngcgvkyhE9YbR293xwNmRaz1xaunZq+dPsQolknKBJL7JhM8N7Ij5DD
ioVIRd+70gHKungYTfCtRI25IQ5qKd4yCHZOYCZSRgzX9WKrYr7sp6Mv4eXfUIG0
vk2NljFYUPKjLynJS0dqHs9W0IEyWmpirdRaRmgpMGRyLtPpj0jC9+wPmLfhG9zp
jBuX51lCdJkK0v9o5F24Ep/bRQ3eyj2F4kpMbuYPXebVY75w8JeWIgdHqu/jD9n/
FCPe5NSSGD/8I4ko+mLPGzMX0oe2idfXUQDDAsK5T6LWzgURTMIz2OON9OcjN3eR
G7Cb2ZelUdjzaajn1mwKs45zVFP+KLRFHtsragXLnOp0wpszL7Q+5jUUE214Ckbc
sBDROxYYQWOmV+sl/rUyfClfq1XvDY7UzPJoLQof5A6B/oicUozdLI0NJOJbuk1J
cCuiaSPbdSzZ8MFk1gWC7WC5o5Ys3YdR6bu2iNnHMT70fYsAkmzCAVV3L8+lkrcK
nB76IZYWEGW6d9eE3IcBJyP/QwGjwK+1YRv1NPksQCATGVTA59gMiEdqEzrGpT0P
MYnufLsMbSvzGTkwE+J6jSAV/34UbTLaC/R/se6pq7zwN4FODf9FYogF5q7YisFK
u+wxqTP12ZiRmXeL2OShVFdrG9QTo7NsmO3Tv2B0n2c7crtEP9R8fWp5H08hniwH
hKy6nhJMwmdT+wN2+kLPf/jIaMvm+nR1qCa0F75iJJBUNeVKH+Y+OvOrFe3ErLs/
7gn38NquR/YorPVbuvjHzxsglsbe4QfziZpZA0GLdao8VbTVNu+tROu1eWNHM5av
sMCe4pbq1MrYUKK9OJvA8WDHHHKmVpASUIh/r6CGi821SxvTpQc1uuWcpB2nSAom
ymZK3NTzNF+EwjcNdb9+v8PenYatt5yYOb8GJYP3Hsy/EOTkBOWQbsIlCg0rFlLh
pSA4CWGCAjqj/IikiVK4inAk9Lqss/E2LFUs+X/viLBx1e7c5KtD2FJ20zmKW50z
Tim6tnJaPWeHdLfrDYoVgcGTrSAUSjXCb+7LPXzgLW9r2w9yHlACrmvP40rR3Eui
x87OrYLnWWFzoruL5nAnFM+vmLCYpOZngsQpgE3i+uFdm7X+4YMmqWaP0P9pIU6B
vIzs07NG8YUdJUuaMUbfIQtP3lD1hEfFlliIjNzLu6qb8PBAesHZkyax7yOX7lj7
6uR3w/jowrYMqhPas1Er3uO6E/yPzMeCnrrEkg0ADn7xCFGdIuY7FNATanG9X8tv
AipabpQiLSX+BmAKp1RgAhCjgj+cCUpdx7a6Vk05y8vxLAGQOHmQl3HONWqWlnNs
0+fzzbGEUfX/f4W4hXv4M/3Ww/PRIlgyP1bnOG9w80LQ2exrN42hhPqf06VNag7x
a74OaWF9oCkktD4BnQ2BhPeDBQKvhODE5sJ7N1hym/zd/3u4B24CKeYDQUe2mAR/
0EfdVUB3G8VA9lpR4eX401wUcHXvVf2fHpzrSDE6ywjQn7AVAaXjlASzN9VEM5nZ
Jn6C5xAJRlAqgup9jtVok6XyLRA7qXpqlNMfQqVTBr8j5DwfISJPtCk1LJT6X7Dl
kbrtgZkRkqsMFVrnsMcqs7yPZthrOjCLO9zdwWS5WNKuvNuyuGw9aGrkP7xTqLaY
XtZ1/0naUhzFmdOX5iByI2WysTNUgfSXqIXsmle19d5nC4cQVuTAWAozUGLGBfGX
WdHEGMdZp4/LkwCKTYqKspvqYWf/cKpkLHyfdAytzk1P0CucQ407DpuptLVkf1fU
XUfCPe9TFVj9Y3Xl7heVQjaZKbZ+Th8tw8fMg8syJp5BbwmH2oU8Vo75HP2wTRNm
XOHU70c9Zs/kCVcTfuTvR0OPddI8qOolJhnNvAKv8bsl+Yc88PLYrzjCxYbEsk1N
aZ8JZzP75xSyVSpznGtnuc9s1vTp1nzhgQwyMjLh6UI8jk6+FXwQ+Ku4e7fKBQmG
TOTWMPNjsuUE8XKq00ZcF7zb7/wkbSW1LVnblYjsGdHHvKH8FpmsltKEilJx91tu
8cgzQ9/4yCKKoIlsX7uRy6sb+MtUf1vNyxFLVQv4qrXgZDzrM4FjYhJ6L1BSphWp
QO/ZmFSviMeVrFvkBM5GEjZ3WyeoP2aZhQShSy9QQkZaO3AGUahZOqJgJw1y5K2t
P50xXr9JZJZSesKYof3xOeUm9hTAiHXlSRHzZhhJ3vDNAFwcGbId3NR2g7EohwbA
BVC92Ko784NuSo3zjBn54HMDdRIvDrcUbi6VOZdRTb867vnaoN+OeVWuRixygZbE
DAqaSzqnCcNt8XD7fxwHLOErcc7x0qRUXKXiz9VebhKzkC+i0kU1wlp4K0RO6/v7
GhHvTTxxe9ZQNv38Y8OhOJINy0SqdnxQ7kL3jDIghEAR9T8pwS61jbZE8i13/oLb
5lMK3OGXk+OvlLse7CGIkMw4RMbuwPAwW6v+0xv5PrK859Dxeg+kCFyN63WzZyH3
3eaCUzoD9hiw/9yaIfbB2gTdCLsYXd10miAQ3GtIqFNK2falGOVzo7S4WLO9X4wZ
NTWgMki8h+z0YYPo/V4DR+HYGkzn2GnNUEOcbfeh3HTnLcfLPlVKRjSsJI/nhgD/
MHc9vaJ2xMyfWU+NX9mAr2/Gpyei9rxmu7j0LiAdwt5Xg1WYDcVkWzoXBbPnUz0G
jMOrY0DX6ZzqKBvd4sW1ct4TU9+qt1c3zeCcVyMqoitcqipq1tEmVZKHSBukGEOw
OcBYFaPtBkUW49y/TG1Fq9a4VlB8HcLozUbNVBAUtiIp3c+lmENFLufDrpQx7eMR
v8zpvS++tq99gWBqiNvIeMi0fWMHl5XFhFO4goPYRK4gjqaHjxwfLNuL9cjNzRHJ
2UqreFUwdbF+JfoIBuGLRnHBihj3lHvi+NbpnrhEw6OgeRrFCjN9fdbS2JZoOV8h
4V+pRx2E5yeG01D4srUPfbyIRvB9SHtaleUjjYnzIuxFMcvjfiEBzJeE3rNWtepd
Rs9QGmiSW6464gAWlAufFcF3TjqObupAFLd+HEI+TAvmCJGlcw1r85HupxmPAfIh
L98jq/e7rNTTSw4O6DiUIC8jhHG1zaI6KVhE5dKfC95NgVrtP1zEll08tRprEwJ0
hbzDdDz+uxwoV4AInTj9fFmWpRSmdsCLimtM3pT4vRua+HPvlrydu7mST48XENxp
pgQxyUbfyif2pypkf2C2W55kXsv9LEoRSYvGapoqw5Fx19DnX5gdL4T7tZh+fQyf
4j/vYIzxYN1Sc/5PlIKCraxSgJEV88zTmK2dl9TTcNkpl5lK7xxFweXvHqMl0Q2C
9HGpR3qeZZloBfpoxCL67al8bXBLRfqrL+bWIsJK/6FRiKA6aiwqWQjV6ddFDbvp
WnLU6iKNF/g8UKK1Z+dHLikF9JvD7KShuTk5pdw2hROYyyCfUMLoLiAz2y2bw9aZ
BZ2DBkhg5juKXkLYT7O0FjjD0nmZryKBO+PUAnR9eN04kcyTivd87cP3i8gtQvEB
1RrtTeJaUFsrel3/o9vilR2wWR3LwLxI6sXu4qEMNdZBElJfVp5mQ3d+t4QO4DNf
DWO/h2gjxHp50zvs33fYi+Nvzju/dUrm28QyWIsjdWmZkX9ZOvfE7fBD+XRCmPkJ
OKltmfcXuypPNCxxUvpw7LBBcXhpVbALsjzWEUbNyYPq5dm2m1DI/4/toy+yBfCF
kguBC7v0TLpzPSznOp8YfYiTVLfarjGSxaYsn0zAD+yEdYpYimdhHBrHj8dfYLqD
bkKj8GbRpe2MTZPk8PnFz5UJO9oFtaZvu1tCi3qghyvXJ3se5rcS/gw/jpZi1VdC
ajUmAO4oJDeVDFq9Dzniplm9Z9JVX1ZMCDDYq2uWKEJgQyztDRUz57V0pjOKsIty
0gbvNuiOflybHqwDQMaN/dv1P+9+y5OQ+Km7rPGgI4B78jh9urG0sF0ImWoRYG7C
KhLFAtstc219elspibOJXEV6ALptv/pbjB48rn5rm5yD7T1EyCPdYhYqpS8xb9+G
YxB7lMkExxIuTmDOzJWqAifVIpbm/ziuTcecKMvMVPq99JPTnCbh8/ses+isMoBs
TBUx85ysWjph0sAkXKqaolD+MMruLh0gB/rZpNRsMmb42HpevI2/Vih+L+wSn46M
SoXnEP/fMHPEjI4Qkl5my7ojLbCwxbBQ5T1ji8faXagzbFQc6gANeuCNo31y7DCr
PFpvtBGMScTjuOx4GnbeYbTZYt+bUIN/tVv04ZkcRp43LQfBAKi2ohhVf9tCxUXR
+0opBW8YMeEeA9ruFRkCP+zhQZeSF6atnv7Q02M18khghgyl4ong2hT4nH12dkos
/fIlkh+HJhtZfuJrorzsJt4/B495ekJb6fnc8x6+OIPt6EDDKal4jdAEMCiwZ7wB
wpmWX6mpqyG3ni5taZNA/NpbZADL+5/eYjoZSyLEHd8=
`protect end_protected