`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 61520 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
S993bpJjwxtMDn0RNN54X1in2kF/jKrxa51VxO9UpT001jXu1v4febRAsl2RYOFr
x/jx/TuNdPenfJpTAlZzJxlRWkenT+TaR4ck8QUUTjWcXcyc/t0zLpX4JRW3ebre
m7pHT/bYjPFvo6mOWIhJBLmGkOnF90/05o5bQAiL+8kbRBWs+mZF+AUJdZJkMExP
Moyomp4VTdZUbHqoryeCYqKEqW5QCCFGvtBb5B+0dKAfClFVxLwGHegyFQML5+9a
SQuSmDz/g/K5yYMTgXbC243DKX+wW2w9bz3yWwoJAAdlrSbw2tI5ZlGzSewOthQW
36Q3Z6r7FtLhAhMl6SZUT5lk4QZc3Ymf3a+Gq5XqbLuiQPuozqeEe5XURl/aC8VP
W4g9yCxiOrFtcE07A0h9ClPvJzfL1OH4jdwHnXLMCIMrwkRAZOdpNDi8roupEK55
LYSqol9EOd0teyVd23oGItbL8cdHA/es7Lb3FBxoxaC1uZNd0befpzcQTc4vkwK7
PM45dIUWGe7qNQ63lqcc9DxevHLwQEiUgzPX0OE/mf+Fnp9NdhQfYnySsTYxXIfj
4HZie9Hb5481+n7Mioi4hC7ULcMI7OOh1YQPp5R4ULhu1TadDVhFWDMPt0zvgBvS
1GnYh/YB556vyTEnUZbl7jAvcSSTzAhhX7AtCFsXNVYbXbWSJvDuxuF16YbUjrbK
fpa3q11T1OPs0nu6zgzqz/HtlopI+b5V/sZt1j1U3h84kT3rFZQUvCmKSiPZBHAm
AkBq38MqlcrOOi20Uv4KKFRWRB9O829EZUIon/leJlByvcPPNtkY+oX+WcviXznw
Y8ew4wo1Ix7rOvuHDRK18h0193sh6R2z/h02UF4ENX8oSVpSCsMzJIDaZhFm1EZm
Rhxp0xiDFWfUaiGhZhF6b6y9PzbEgtwn8M3JhjMCQAnryCt42qUBX6edLnLHCpIj
X9q7pZJBFe0knI0jh/SDD9/gIzktw6uefHRSAE6sLVnoHrDGuorHuPOIEUmDS20T
88wbp1BlKnpVXIQOhRFSpIQX+YeZZOLZCf5lcsdK6qgmsXjmMwFLU3SC8aDFpa9h
s3RkYPH5EhzmP6RCgfMM0mLgLzx0xPC/4rQg1dxhF6VU7616dNcOvN5B/3mqK0Br
gp8S5XaJnPnpmRgp4ubcj85VEFI7dOECeErrTfjTXBhmwf2G7+2LKXaXpecBqxB8
jZwjrK7XhK2SbRHiYUea83D4X+SaCqb9zIQWKK5NWetysIw2ylYkK6DSRLVfiqEG
k4+BasFFjZ7D+beW2gs1rZJsZJ33+KJrMjokOPqLlA68lHYy83ElTcliQzPJ8rJy
Byr/bfw5uznCd6iPi8pGiXWSiNBrCbpFIEEuwjQ6a638iWs3N30GTOuWM2TzvzYl
5EAFOxNYbKIVEVDAvyuiKGHCvoD3xPQNvbARAKD6XKZuJ7h+9NH9m6cvfEM3O9cF
bCDzazVpJxj5L0r90jZ90/C8FMimzZIEhJwVi1zwbxSe78IMA/xubDK/UV/sji4j
HI7QuEqkhFVlwI7uNAL1CBd0iVqAVtqMHN1TOqeshwHynq4mgqo1in5uCFENXQLv
syTTSzqU9XPk/rXID09eoajCMr/ydAsDzMy8WiNI89bVlDD1Q7CpO3UaipKIYaal
i/XvmVE4EMo5ovr4H92IGv9nr74D3jJu8AzraNNgiT0Bn+6f7th2BwCwn9wPx4NW
fNL5Cy+3IVFeBlljvUOyiV8FsnMVCcA+sLMA1NjhnASd0e90WK1HqWYFhoVKMoNp
F+PciXPDc5l7xqqhND5fryPc4Q19Bm2rwd7FOFIHcPQMy9/oPlYEPZY5wUCFVzN7
14tXO+VgZIbDRf0f5bQyMdxUXIHQwg9bWeoW5V7iZkUh6VonCZ9pc+yO0q7hBbxA
nkr39NAn22Jsy3AGhqR6HXYgLVsjF212fKPmg8P10NLiYm0hMzBzGvqnFJVt4x3X
fBeGpD6Ndl+TRFQvl4TQzNbSNax4gbkegAAQVK89+NH2UwysP26OzdZoOluo3fsJ
EHImssMGYgBN+VKbuA6sowiMg0TcK8fGXcqcWEH6vURH9pYVWhzb4SCDTSgy2npH
YWMGc59SxTey/IHHvJcQ5d9uG6kQDp/38LVMJZReIx2rAS/MAbFykUrQ2EukzzLT
/6Y+EjMsEojiXm3cEVJs75zMRQQzKHlDxWVnqWcoxQotn2UAhE4iw+g8VuVfYjlb
1ZqxpdCsTUUS5qecKXv7bsNw8DaLGa8BkLAf8fvkEAhattjGtExXee5Rih8ERGBW
W/VSCwLGoYZ+2HwkjIlww2jeJw/vIjZja52vPdG1hjfu1KJl2q+SkdgUzqgwMQgE
WRW9tv/FAbxfxqOUKUO8kocyr2NGYx2hAdKZOWvZFXk3pwSXoQEZBiuITukop1Pd
ulgOoQdySSmyunKE2BIN/S3mOSqzCbUINkFgzYYnsfcsL0rK3F9MsrYbbyRJLrwr
16h0ij2i/TBLhNCSsDrNeylKGX6cDz6TKHQlx5numgpqsdm7ftWlAapcwskD0XcU
/hO2FTSnlv9gWChfWwXEvMTaP/eO0x2dtLglSVlvk360wbtO9ZVJyvqDflYLBn+e
a9LTN+RY6Ah15GNCojNNVxzUQzQcHUzrzbddAFbM1Ol4HAF6IXSg8W+u50P6qlV8
78/ZnpZdUm8hXe666XrsuqIBVJOo/0P4dPsen6mQrtbVdjOVUNfhwVsl0Ov4UoZb
f4dIquFAufY9pLTOvD3RwtmiWaIX0qtgGnICMnb9Wb3r9PRZ8XaJYOCY+aIfFV6L
MD6fWvUKVcwUcWz6dODW5fIghUKV0gcABIxg0lGLsCHPVVc4+2bmR1M3u6dDATyq
uneZebIdKBcpom87im3Dk3U/nbn1dpzLe35yRpnxDqPH2VewmVvaFXVrUEaIm9Wa
47rbM9fFiiyXQ/DftoWWgp8+sQUcxvfQyNBj3zcDZYg6E4S05V008y9Xar6LfCCg
DJStQpS30OS3sRulV58cOSSeHSbduTj2DaClxqsetgCsx50S84Xjn+oa6lvUNQkt
cCciIPU/XZUGJpZDdEgCNfzdgVbLWJV7hnCfMGX3g9gtn+rPF3wyWwJ+73b5LyKF
Yzj9+SS2qZR+xN6ALRsqyIQomD+fZmuKCvjaRp2YHy4izufJWJZQTdPcFkCCAEEM
4i0MJLTN3wDBq8hwwoGomy+5q9Tz7pwD+2rDc6falmR5UlKw+se6t2fpDc4OKsMM
SnF77a8x+3CTrpx+ASWe8h7ZAdDRF4MnGLWiEMJGcfy4ghnweuBTc47AKWZMsVcM
PimA6uFi0OFzu3Grz/DmBIZRfvSTQ+6byM4UVHCKNjj0U4U3H5Tqjk3FZgosC7ar
BgKV0hTy+2ZEqBjhmkZUT9vvDMsq3t8FozZTAoAqDW6WIixRkBi0aPWiCnjO0M8t
j2eNAwj4NxoULEicuIfUkd7K9OTgzy696nSu0fO0mjOdmDLwKLO0lFxB2u5bacrZ
TDo0kTdUX1Q6cc9Y8sY2L2RyiWJ2rN82Na3Lp+86p0S1bfJKL9R0lfcoa+DShK6f
N5rG4eZpgK7oriJtwAkf2gSSi4eElAmtzD0MsTYhcEswK689onBqPzryL9rE+O9I
pw7qALn6qDAI9U3/bQyCYLjBxfHDNO36x4xkslZ3gdvrO16cdAXW5XZTk9/+ERK2
xSfMpm48kI6nc6PLTw+lJEmHnHdswZjUxrqZiWB1E9DHb0LUC0Tp4hFl8Vd22+2j
jR7/zDfNd1tyACZJKbkTD9FQOEVbAeSwLpG3Io//wWF6KxBDd4sPMIjH0l07aZfh
aIzCmNw6snnEZTcQrho1ZDRqhJcUFyJ5QBNG8izdQ2wG9Zrv+EEG7bcuynzMu+i6
UTbgA2pq15JEGyms7aSbQcCCbwr8V8Q6EiaqaZng4hcQ/aIgvQxxRfsEKAK5FFlN
+ElvDKejfAUJFXiWdSnuXb4gAJuPP3pvbEiT0sG4PQ5HmpOzTkfMbDLux7agtWEF
Amu7L33bVLufkLSW/kBdj4iA0/wdUQVcsp2Z5xk4YceBrQLknOl6VFtdIyfQ7KAx
nrGFu4FqJofgLBTBmDGgkrhCN3mZDYNqTua7YTpZtBl/QDHCHBMtat4GOBJ0LURU
heEIrhh3gvw55WoWTwgVgUEkjmlRUV1M9sb8SUQT1tx48PVW8c8NGGw3WCsC1S/8
FDvhIIMpIRozyAWsuofol8/okzb4cvMAvggccNEyINUPd4I7RBB9pHCPU4ooJ8Js
QdrTbpK5LG1HoIPDT2mjSJmIuxJMUuSoutf5s0UAflonqQWpsjGCm2N4OzKi+wSV
nPfl+pyJcEYWNbnw5tFzdGxWS4gAhbl510+Y074zuKWfeWMxsBMbf/7451ZWPQLL
5hwti5MzCDUMyMpIYsOHqIB2JvVMpg9tze5yVfv+V+OJm0b8xNi4XtXyc71KO0NH
VZ4MDLq4JtoXeM24WsBBr5bZIFYBRr4y9fcB7HN5tNaUJ+3SR1TEuqMQrHl5G0bR
w2EvEqLYhPzTPdpiDprlViMA3Yxe9pdNmy2WUirRbFe2fQSnee8QtJGMVU6bb342
e679iJQrYB1mWIxQgbhLtnyIJ7oP6jfRahzkHJZDtJLIlcHLjzt5+HmNHQLTC0Tx
xKUKgRmetbChYcdmEIcyfzGT38jN4HhEP4KFOTQTP2BA3xDCCE39Ot6TMf53dRp9
o6roaPw7vDEDEkDkbd8Q5lOqTfP03zKgIjRBZm8WpLM3fyxUMX8vonflSdC+x+D0
/R98dzZT1Jcpi1c6/YShmsuMVEN0tmNJMQtDrhbUI7BFbHHS930VXeug1kD5E7S0
lSHwKA4/8vvGdIz3WwbI/esfgGpU3nDXCMEHkg6sAF2y4T69676fiuk43m464Q8h
q/mi216D/06+HfBqk5jUp+1hRPoB9FJ2U2q3GVDZ0AnPButmpIy4grbNy2sKzaeq
WbYSrNCQmo75DwoxjiZCxQa4xDO5BVxLsKWyFN8kmp8nDtzX6gvpXdp2wU1vkefN
ipgvLDNYGA/BTIHWSV5lulbzjZzQ47jJ4+8iFj0Vrttwa7/hB3m8CoMWxYB5FIbo
gxG33nQmyD1zhqTee5kJpN32uZDjUf1ogaknuUyL46biDzi15GNL/PTfBtjYeBsu
Fn5F74h4P1HyYow7E6WkBnVN9aAqjmYyiLAF4jmH5BIgU6EutxlLHpgw8kizLzGc
atIjInm58VLByoigtqUBxOgbUPCUtBDLBCrduNlf5+fNA9qcTrP2abB0FAHCbt4c
ojpDyINbhrKWT9lXsSBppXoH88mUz+flQywMdLQNnhIyZoBOR5+J3Bz+I89jCNRf
cq4h2/8rmuBmty8088xaYoPF9YwLuHGLxVY82mSeSWhxXz7hEntJU6Apk4ZxZGcN
+86FDOm9FbEu/yTJ2D5EHXeZLAwrAZZ00XhDcDSSbz5ei6o4pbSsp/CqhaCARW0g
JRyjOM+fiPx7NmpEm2hh5QuqX5XfE9A8G+K0x/bJCSOfW9ymZay0ci4nDuRxkyuR
XKhxj/yHWRX1sIYHypAx0dTC77cVo+my+Sf4AQpjbelmZ6jHZ6KOv3gjAAXhxjrb
ab3kn5Vvy1odUI82oX0QqOczVsZoSAPJa17acN/QW2BTvPvwJSj2n3kfWduPn2mK
kbOrrZ78V3wjIFTam2omK7sSO1U1WjfiUfPUZ4YlIJuHcoHQV1a43W1Qpcc+vhU3
mfK4DSM2G30z4o7viuVeNK+F0vkAyw7TrI1fTA2gacVpU2sEbr6fFqTMbg0V9pUt
gTcI2tB39tbwtIq9IoKnoZrZchvo+ynWFoCMBYGxFzMTHgKNn3l/QX26ugoJJIZ1
dde32aoXhERTUzeFVZpvr4TF1FHGqcJ4dx3cwpk4/qhAh+oA1qduXqyAxtfvHKbP
vd3vMBAJq4D3ykttRuvJeE6Lw/JqdHvstckyKHfLfoZz6WN14WIaqY2SyNpI2vng
VFvENWV5lpm3U1GVYvfQe0k1Hxvsi6ycTpkuxpdkDQ+DpgISuP7TopdJ9VlChzye
pGiaaGUeePbF7BKgjYvymYOkxEUN6asbeRc0ROg/jlbIxX2LylJHqX7XQmQMsnsM
5fko1rGRzQEA08W4NSGcBLk3aCYSP3Lu2x0wwOy2WS6x5dxVJnzdx29u2CJ2FuK6
lUrUF9Sx1Y6pYx4O+n7XBsJmCFfvxlesXeFnxNJHp2R2UeoFflLVUUKpgbACKU4m
pM1bpELaBNODDn1WRfO5lRxLqNUXEd/E3qvWRVNIXd2czb9WN8O0Ch4lJrMd0vhF
KPu7hKru0yHDwG+Gz5bmltAFsXYlYXGG6446rNXS/Vots/5HEWcwNdwcqMXyuDGE
eJ9lBWSayXx8aM+n4D12PoOjei/hH3m52uUEUhPSVtf/X7OWgoS1k0wXR5BmELrc
eU9cllU0LI0cbotYyAysVJvO9A76QebQbcUHuhmsB7IH6Hm5278yFyV4fCxU0jaC
PRaKmVwkT6ldNBisI0z0Q+N8qBg6bceKHADxTc/stXEp6XSUb1coY+K7SX9z+EIM
SMTAGAMm8tJr8DoHlINe8jxY2Pi0KdS5g3BB0kj2kZ8Rsae+AANiGdM0UtjTJIfr
i54ZDkDw0RSpmO8tFCsU6QTVQCwI2YVyuPdTYOsYE6A+PvHFiWa9xE3bAmTHMeP6
+eWL/YFiTAl599g4Tt2xrNq0q8lbMAssBBPksQztq/HVqt4u4YWmGGsUY1IPcUNa
GOPj0yrMaUxKBsbQuAqS4uoA0YRfr2DT3MvtK1KqVy8paSGWksRb7K3U1EHpIYS4
nfyfYlxHCPA9DIydHYpy9PppFmklFSFPvSgCFG/VM1l0bSQO6qPW66c87Q6pGHn3
/dYs2OEc6HnHzEeNkzXbgi2wJ9/EDx7XfIo+ZYNQd7S+lvzLXPBrkV/LjQEHgPCz
9RGg+djhB3vzpPD73hzbToThqbFJwKxNRd0s7hT0Zu8V3pPC0sQffJ96a67eT/2c
sF1YAOQAUfcX3Fi3hF2nWW+9h3o/pfGqMWCv9KgO+KVWWVvcShosuXAJcmoJlxoM
qx5c5YzthJHYvAcRawNFnjgNqBdkcJv54eyed8c8YcgSEASQAaXyNzYx40OvnG7L
Q1UmcLmU/1XE6brZ2plzlS7bMIsx+J1UUH9VQmpYavPtubPdvplIMuvxGSA1UBMW
XrD6Z2mieUZViLQWGdQXFGB1G+oE9tbG0EvPUt6pUu7wOnqRaOeiBEf1Uwd5v1Wd
DBMCL0oiT+rShDQ1WwjJKylEjamgiUuyQYsdaOB8Jiy48s1YLDsyBINOJt3rogBk
V8ym56WQPCvd1KgDV/fAcz0FCAg87ymiIf02PzWhVdqpw45vWX/KXVx9WtTkrFxd
GCc0Z8FTVajrVR4WRQve9ah4ZxFAerMvXf7ndZOO4oOVnMa3SeCTWd77GGMw5fff
R/kF0OtLhINlbDlaUGdY5fotJAY9d4T7SnkbxadF3stxhglhsnwc++GTIpGEtZwi
i/unROYLXjQ0lSwUIJLU8pzdLc4if6M+k8bDM979zTXUVfzumYaJchMNFOVhuaD+
VkIY8v0/T+QphKdktMbidiuuQsLCvtEJVeUX+/aYPpT9QYNbZV58yVRSrXJjOABO
yI1Tr+T+bZgXDwUjnhqto8r5UQgjN3XLPqN7yxzdsHIV0HlR7Eg1O7y2SrdxfYyy
JMCcM0DZje5uGACUvXxXLnbfIp+RXRTM42VRAR1h+1lnw0lSJdlxKShf4DyYIKlY
XLQSp9RX/xYLnKISqd+1qMNMk8kiZHAvxDY3EIL4BTh2EBRVnaRArfeShcPbsCHx
5Z5vYPQ8hC1InnhjxpKi3pOmqN/RMHFFEccEsU0K9OKPSF87SoAsjOryNFUnwaid
nM3401hjyAKehFdtz08vvmNOz56JQYyalbje6hu1OSe4Gn456hGyttlRnI1UqiDn
SYxE/fbXuIBrXM67QlYRuYkY0do6qqbJjoR8HyBD8l+JKXTsWMoiO9wWhJ3pt4fW
4K7DAP/RfgDYNWMNb5YS66QxdPfK6xE9YZmI7QgyCYbG8j7vU1RRIulQcMwZ5HQG
PPmIOHIsPn6k4IquTFu2EuQhTbx91C1CbtB7aT1V/PDuC1DqONjcErrxFLsaJXBb
nsahHuMJUqIF3GYUhfwceQXzv67qTYQJU7Izk58jtqD63D8D1nQAXmCvNIUzug8n
pQKe/7ewDS6fw0hKQW80+v2WIy4nQrfLX55fvmjZ6w4d7O746WPKAnTwVNr64IiK
QztM5v/84tqcBCemCSzc4TwHPKK59Oi/yx6OwuQi8dP8WLiv1aDsYkPQ9ffH/0CG
G6oBSy8JtnDxMtckv51VE0vRp+XbaK47F12YAEk8keEz/EPrJi9MBTCyVQ+U2vLN
Yakuok8+rsyILF098W2OiI4n/4j4sQOlbA30yspUoyJDBkRkBnHPAyaF2siis5BW
f+wczLadM9sFiQhARp0XVqTcG1cRPNUHSeQYzYItrZr5FxQaFHzIJbiTuef54+p6
SgdkSWtxviK4pQUWs6adjWiGAnvZzgbKNWyn3ASCMAI+R85+ji8wpbZhe567UReG
RlG8Ugmc+imz9rsOMs2AkxYRzczsoWAL4H2CpTQLFbOBUUKr8PKgnzjresSag1d1
JOsIiExDXe2ab9ydHq4RlXFe7WtMVjgmT0FSKy0VM2V0bt+NwRbREHPdAlqwf+qH
fXfp7RaCtZY+9O6sSb+O/IikYC/y9dbdizXV+NqZ+LO56qk9mH2w2OhvaVlkbCJo
MytD4D63P6q28QSGDLS/Nt1fyVoruIlusrsZBm77VAhMUBgZFXSpNrY8UwQKP/vG
U3sLVZp85CFWL/OUhgWpp3StUv95xwD/ulTx0Cuv1YFR3zhDw0YQ1zfzRhzhbuSz
Dpele24lZ9fzLkKPWL3bgxewm5eNZGEBEUh7HAApYPYi1yMHIksnOMW5pjaig9Wr
FLK5J/oM+pgrLy5FUPiaY+E9ko8/YMWAVb9SMaz7icEMhOW0Hf7jSGsTW9e0BSqV
UOmVRO1lcipxVCmdg9IGflpuWxarH8PEUsKzPYLgbskTSuyc8K+Aivwc3XyA5bIO
voK+02DmaceEix6JkwTS0mBHrfrS23HK00TkvQaaWd9detZjZlNZYNlvVQ6oWjDO
PRowpEqhS5zLkjIBFsbVYY/ZRJfOOAmQZHKescq/tdbD8cJ3jK9IRaPuY5br1FXo
NBaOtGnWglBEnyNl1R9SKwpuzOYE3rm8d8nooEFzX4i+pt4IFQyw7CT9H0vc8AVA
2jMgFUFeZHE81SZpiNnBU75Fclh0tgmbG20NAFg+lYn0KHMmg6ii/lMM6z1xn2Mb
xe0p+dwAoUCZqWZRg58bXR9wDcqyLjOc6iPpeBk6n8e2YyTxJ51PK5GpjgJ22zLH
PLKH4nGDR9Zowgx4NIFKZ+6qxmNnEWtfdgGLZDnblwzoePCBqGPPcgae7hVWXpk5
iq0zX0mVtbmW7v5wm+ClYb+V7Y2iidwiPac+j+MEma503d5JMz2LsCKPeLz3aNSH
QUw7aamrfevywnQHPC0P8yKMhy2os5bf4F85lcMAuwrybsQCwrvgiMKLK234W9Uk
Jb/zSwsH4Sd173KG56+nDg+EiJbnbsN42jzObkNSQn367rutrGhJeghBxKPLK+N+
jPjJ4GYG1XhENwnqRNreSYjIhzHel4fzx/jU/TWf0fOad6rE/EKw3+Jl4fN5CszD
4H4Yg4Dlc9lX8LIat1PLOpmTRr1g2KxhnfHVMfbS+WrATrxijNqz0fqL2D8YSAX7
r6BxsX+JcUIXhf+2O3HDR/7XVvvXl9xjlA2zdh8LtIMkyJCRxCYqH7jPQ4t/mvJT
gPb0QWWGyJVaxoaZDIp00k5LbFHyZ5dTq8IghjV6hZm3a2w5dU9IBkaEQH8gSDY9
TtsBbpPgj/WKdn3/zGusk4xcfdo6pKuq1JswKKLSro8YUcyz5BV+j6iFDbJGlToj
HAR6BweexGXURTmLPfZyk/PR/Gto3FK/KcN/76zQojzv7v8lGZGmsJIGtE5nzmeH
3H9XW40mZcpeOWLMz+pFUhtzFiR2KPtyzAjnOzec4ltsgSfmzHHga18CMtAmT1OU
pVX6nehYkXpw2m5QD6FpO6rPIxMccOvQ9lKS+seUDD9ElKitDsdzq9PHi6YyaUjo
hrRxUUnIPxhNW+D9J8bCGzwCvajoxJ1g4uH9ikvzx4jiTXzyS77QlDhbOYiyliby
ROez4apKyDdpY1OE8N3YXNyBisg0gWLqXR7oWgxpZZHIS2LmvNG/+foi8oZrra1U
b8SDHBvPegzwkIiSflVa+H0TjqG39bFKViuxwVbu9JftEWeCGL5Mjf8JBiW6Xe31
yfsual92CZhl/gxGo3Lo0iwGkixhB8/Onvo0Oyg7opI1YrApbroll4+HaOnXNUtP
mAwAGf6HII3/acbO5fSrDh1sTO2+NLkY7hoZRrUnIfKUeqv/gQRD8+XJOepaG87q
7plB4aH0Z3KYCEy3FIwQ2KrUj5qFYdI5UOUvAd8DaLm9h9SL3VDHYsZdGqj8zHXM
Vk5mqMeemmOM4gHRLMUKGuSa7IEGPz/Fh2dNbdaYmXmI4vFNIj2vc4EImM0MR7MK
Owh4CRLhucuI4uQgF4SPT1rxAS7I77kJaUOJZ/ioYow/T46+LHQWO1Yk/ApXjz7w
IciupOgocvIpPJIBf98s3BJLh1bbzGZUp5kgBS7Ao1AwEWe1su6iY+OPTrC8zUp6
QOEwl84wr+0kvnTzHWWegMy2prmoidpyPtAaeKMfPEDm6qEN4SIFPgrI5FE5hzKi
yTYG74CgG86+blcjBPIQsp0zY6Kp3t5JnbOVKesMbs13p8z2405RwmUXP/zm6vKn
ld57xm+0YMvQ4uumTyPzd0LcIPJRpyiRicptb/WdXl3zuJCGUXfmVuOBhjs3USRC
nqNt0xK0e0TakV+YtsUYmh94AjDhJUXWRtgJalio7NgBvix2n//s6K4l1pCsjGpE
gEFG2e6Mo7Q+ywfl1yfWpcHWde72Xs3ssmxdcE7Ya8oVnVLtq/AtoOUtn3ZrGb8q
YaCxJ9hnJEVXBYwPInXSnwvRc2yOICgcdAy0KvN1VgASqD+EZqLk+j0KOQoNgLsN
WKmQr6mWJSZuTRDXZow/Zwz8r5eVUdlfb3TrZTCTYIi91Wi/Lm/7VBlhJihXTXVQ
s6vBuuhG9iUPu6JFOi7Wiw1YCHtA4rzSnoM+cAJgZF8bXp3rJ7Rkd5hyCfvPqytA
ngLTEkQ74Zat6Z7yIikLu+lgwsShHfqE/Pf4UO8xtoqvfKOa7QJpX2rVm156FsIr
b8z+ap6pSYCFXJ4yeF8yMOaGNmDsiESO6eKMsxFEdnjUBc9//nSlUHt/w6fveJ7Q
FrLsuaYK7CV6mKSjKu26j8fm4GGNyRZC8R1uG3VObKUKX4JT4iKewSXIwu2ec2FB
yudVPoiACSetHsiUft6av+ZllItdLUpPZm2AMcjoVJ/Jj5hBX8D/hcaavqEvAtd7
59c2ihA6knKbjvXtBBuwONHDbApSIg9lS0AM26gBNaGzpm+7Vyz6u5SGAJ/i9+zs
zwpUjZWvDoDlat1W4JIHFES31xelHE3qfrw1tri6fT8E4K3G3O2/efmL/dVbm0EU
5LIVFMDfSCGSxMOJv5YxtyCde95kqayjQdaR9/Pv94vMZ8aqr3ZN+/LS+/Dc586W
ihuV0tInsPXF2unKhG9Yaeo8ZptLmz6DHLM7GgN9Gth/ayQazH27ToEwn7XncH9K
MHN/3V2jMEGNijTg6MtRReFS9C6M/4/REXN6dF9S5kINGyGgmbqCKPZ7Y281Skxp
dZUWIAdUbIssFdoU6tI+VR96oceylygRhSH4vgfOuKtcHAkHJduExrBMRGdEL7dG
pF6marAx7+Zhueqb6booHNkGvO1I767o/LBB+lRUySKmSQplVxfLAEY3tmvX9EsT
1ARzBZOjsWIUwTqEUtP5j6qUGmymtu8JoS1iwJ5sY1kRbFTOO21N/95570wcmiOl
sHrtkCShZaIKps2GFlR5YZBGFWXZx92nA16GnfxbzL5zZ9JEH3P7a3qamTO6zDnV
27VKW5In9XgYh41Q3q0WAq2SXah67sP1Ui+UVXdcqcvlbjcQYZfjJD/QVGW5zT2P
Rgg+J7G771S62VwF38TU/5Yk7emU/r0z0aSaHx7KgYp4qteAl4vyy9l82pI8UU3/
YsagYE8xa6fu1obL8PqRyd7AH6ytxEgvXG60kBz1L1mSsZDZuBCJB6zcioNDJmM5
VEaqPxz9GSJ+LHMrPJpLK+NNX/H/uIZDpN6W+ZICe8GQT5hDqqzBZybMirpX9Psd
m7ES7DnvJUTXy3UDeWlHkovDmgVXDPtT7gENOkvyRWJjwEmluZWsah5d2EPAYadd
13/TeYxgBiB/18yenWNu+rqxjEryZ4Lo9eMjb0jRo15OAGxlrvCrWUMWVAqsS3aV
MglIarnXRCNn4aanAqZOMcJAikFZnkFeXyx0ISxsbpQFhi1p5EGbGEyk+aklcjO9
K5OhZH/3xbbt1DK1dxqhpywkzqfB4CjOGnX3/Bp+l0iQNsIAQXJAUtLTrmSkhYfH
uPBVKOADwDCSKXdQLM28eEl+5SOS/EFBse/No4ZP6sSZ1RJZ/PLrcUzZ0S5YoT+l
reUsRSMqGlQ5qCc/O1EPz8F4Zjh14Dv7gR3tcr3PTNwQrvuV/9VF1MYSUshcooWJ
2YB2j/4m1rbwZrJDBJRuNcRJb382co9xALzuwN0Nsp4xHH/8hTxUP4ss31bnuUoP
3v68xgDzxja2lGqL9ZVdigFMKlql5jXrodhKkK20ewa6uIuEx69yMqknrIQziIg1
Q26hoWxMLBDb8wAszRRrSQ+YTVj8f7tCvOwBGlzK+N3qTHQe1h7prqqucBduOpLb
YVcMUg+b5oULTX2R5CFQOvP0xltnak/eSswrL2+zdjOatlfwSEr88iqDt4zmk4DE
lMJN8t3OvkNV26zwJggeSP1KqJTKKyEP8NpveSm05MMZ/KpWFRYetCxnxW596shc
g7f5pd53U87TajEGeZDZPI8OeqMdJ+ox3X6hFDXppkHGfEK+jQF/ERq8OUvMeTLX
Oo88+PbkZOlmoaCm7hYWnaOHM3yM4KJiQSsJSslCxZErBVr5AIU0gtpvz+rbfdjw
Qqme6v0OcNS5+VnUHn6TQtDPT5aBvA8BGnmkOIM/oA3qISO7m4ObSm1MKTjVC2q8
g7nq+pwc9gjSxtyEN+uueLmsiQslbNgD+/GIJnp2288406dtyWR2xMgBQZNway4z
qmyWASSOPmsMshmnmg+fEW1DqB+yUS4tddPLJtr1ihx1MwaZCai9Px/1VLLMUw9Y
ADNITKpy2KT1VTbnL9ijB9Kqh6+37Bax4DIll5JiJv3Km9RBjC9y8KofrvoEMvaR
rQB8bJWM9V60dWhlN3RMSP4l/cftXTFIFNdUvo24s5t89T+71XAfy3hqYt8XQ9SH
B0yLFBP3TiQIu+geFbBjZzXcYVcNeKiAh8+k76d6iJv2+wTUCt9L1PAmWAqMcf76
Cf6zJKA0bohN9mlXKrFeZenY7AcyMFKZ+p1rvxV0JbfHBGouXYQvGQJMFtINdvKu
EM/Vvdy2a1uHZNdbVBRg8PbUrVw/gQbU8KQzJmN1D/QrurljoasP9Jf1smlheR4k
Md80RVUMjK3/uzFmp6XMpiAy3A/q2giHZskK4Ua8L1+u6E2/mj/yKwRHnkdhtJxj
8Dg/T14fkVZOQumQJC8PCntCRxrJnp7Hw1VOt3SsCFjlAnEQnJUqUEOP1O2iWVkb
DGYYuC8A4R9d8PtUAW63fwC5f7ZxGqCDcM90ByxxTKMw69aOvShit3mh35Q77S2S
FCdPjogEWEMt83swxChRuX6vIvb6oaH+qxgqYNHXezoyrstVdnHtfBj5KFfqUsr7
EyWYTpRGLC+uvhWRm4BoujNsIdn26SSSC9uFvaT0erRXyGJZpwEKXDW+j5KAnjDv
wYayqAjUWTDASR6blvMvp82NQpPvNUDsgMhbRrAeG0nSo7ei/TLBtZ5DICeXCl2p
wzlBGHBQRdkItebfCOK7kdlu3dPYvXz2MPpC/rGwCM3TBduGqJnsolCaVbl8L+2Y
ON0zit2QkpA9JhsAZEvRS6jnnc/idPp+iVmsMYEWBI5//J63P7d+QURfX8rbBlCP
JxX2Kpa+puXWcr2/g3nL2uulLehSIP80aoHXqqhQn1dLOsT+xHnyB4psQTJkIZSA
7lgU5bUePIQcvDDiKBYH4paPXPx3TdUGJLhNCnA8RfL4cLVo+/27mZ51PrD1L/9H
CRG8Hcv8Ms6hAY3v6ZCkoeNg/2v5CtHRPepMQM/r3RcFjAIeQOSWgYAMFrgT4ra+
ItIdEyTt+rSWx5zZu0uI1iU3Ss35CsoehfthihKlT6VtefWx3kq4+kQtS0mj45ZS
fJIMjuFvRsuYsonCYn4V06SS4ZnfWTGwJ8LWoM0otJDnFHy8o728R1BX4MmCvM6d
cv+BayWhMh9FqkA+8Y1e2N9qRGOTiaKBTWHGhIs2/fOdckaLKqrrX1l7Wq1QJnut
etuzxFs6C6pifetDhGmprwSeoBJXcmtQc4ZPAghY7qM649XGSnTgnG+tQ3GGv5GB
xtlOmvu4iy8iyzKBxZ+uplYsvVkg6MUpxq63gH6rO2BbYHkeZgPjlRW3MyCx5HgX
LYAck6gy2eu9dq5IKab4ZotKSwLbUGlyxqg8FYW8bUh6xdlEaae4xbhX+pVsLjnj
Sy5WAWXVpoaYCqyh8o6jn/r3i1XettWwwvg6k0wewPIjcYBjujGIUark1ZmK39WE
LWo0WqJcw+G+vdhBfKoJEenMVmkDx8KJJjCjMRXFIG4aAMSbAmZG0xoAwE8oU1jN
HgnRF+X6/+f4AaKGjhyWcykeawlHkIX+GlEMPnDocD6drRXrz/ID0t5nqKSqxZQD
srOs+5AAOkKDhbT1VYr9m8gar2ADLg/7B0Ki7CVSYWnOg8++bO1TLCVxltz1+ypB
6JV5TAPoXu3xqArpl4JDHcXW7KoVx/++KBpv4iqlVPlUURHcR5xKsz+1VY5wzjFs
KMLM0chi9sGlqGiJlaFUJ8B8vCKVAQaxUByQTXO/cI0uktuv77M2PP9kr5VMzPIC
8dlfQpTyaT/PdCGfyliu6eNaD3ayUcLoC+mNTU+ZTxpwAURsfiGdE405pIkWN6dZ
Oygpc4Y+KiQCxWaFjDjIlzMsfWQq+ie9HMDPz1C9y1dadSXjMT2WBZxvxa60VWyD
kUxTTNogEW6rJm0Y83wAHSsrq4yDpSJfO8HU88IJaRirCtiwYS1sAmShSG3ydC/6
v+QTZ5FHfSZxv3Etr9uNWEvrRcM38mEABBy0y4FRAqgbBIC8aV17m5z3cp+dHWN6
HjAI52te9GFCJPreeYi78royr7nMRucwFEAkKv88YULnZlbJiAuTO8xfviwmWh4K
yWyyiIMKVxCDKfQuvEUW0/6/4EEh7vD1LGreGPW+XHnmEQSSevXKuQma5tY2N66P
MqVV6bOTbsLp6RCtRmTRG08APQJq7EYPGgqonC+7qcSaJD3L/UeY9u2zayejHCS0
EDXUJKANOvgYzvTIoqjDpJhvawUSKbp3yzIuVhbAtR1D7QYUwKqTZ1g7UsI+v3dK
Dj1lJRAR1pGgcnrgvbp6vpQ8+Fve9Yly+wQXqaJv/KHaf5xprD1ibXbvOo2Wj/73
BTA07ixr4qzWEGIxXWTzMXEpsXe1nBYKwFEgICcOg2dwkSKez+nRMMeikUTlFMOM
XTs4B6GZeNB7boH+yYLTm2Y0i1/WfHD+dVH1hsdKNqzXo8FFUuAXZDT9Va2af9lX
2vAoWa/xeI+NFAPmd4gaIl32QyRCjdm+pQWMnWbfVSeEUMLVWQQrqtKR7orMfsVY
yPxaIxqPfFFWRJ25+bvgspLNnMbqWf1kQVQj9ggJZcaxCXfk49PAFnJm8tUk0Psa
AxPdHx89nlwIZ5JWk0vBkj0f5poPhFOdDmc+I1OPDZ0xjC+kFFyf2P5ancHdzRN/
p96oPD1T1MX+zHhTpHlCfEuH+r9cJGhc6HBzyeNB4yCuKgbo9ZPQq43XtqfIa97J
gH5g36EhYnQ5+c+fxuFj4kyaQKBV5D8xJh4t8Hl5aj1qvBeEr0kUq1Bsx7r0drfV
RaexUPh7ObDrJ1akCKCbET48ny6yBVNDA+Hbda3FrwOOtCZKIRRGaX2CIfcFfCMS
BnXm56wZFdOOhohKqYFQpzQephZykixDUiDC03Hb3d3exx2+RRklmIiJALvfv79Y
HDTadfBuWD05ErZPT+P70x0QeEJUk2vAbxX6PdvoP3Zo8PkQINrEnKtOF8vJyaWZ
ZBMXlishlK7MWvX3ADDW5me+Zma/5BzDY6iUw0bTTcA2wZcVrjLjaKHmj9EMFTak
wJYx1M5Er4Pii1M+N88RxplTeC3dlbmv6+qgF2ji9P10P0nxyWTpWv9PUA6HBZNA
iYB3WefkPZAT2SmFzOox2TPrHbj6ibJ3q57RyaqGKyVXRfIw755RfNabdxkJNN0L
veG34qt4m/D+xV6tqtvR4nk6der92T6jXUO02Pq4qG9DOePPAmz2DJ22rcos99ll
rrlyMBePuUDe0dK4Z0cQLXV8OO8Yqyvr6PJ4KHxkZujE3Gx7hvScbV0jsnQ1oR/c
wcbSEzkvGj0UIjdHpCwYzxQ6G+1z44Jsj3hh7ATfJrGkAn/rDGLCd2lWZnjDbJBd
oTAnDzyOwwY4cJdIMPqc8tkYlwLe5Ep3GPgZ+H5UQcGn7CpjvWXyNmuLkOXhXwPz
7XbKHb1XZ7jprocimqL6IMJt4/ASt7uJi/mN1nAAGWnm8PYlBwIDxVOSkl70tK6t
Vuyig/79pch6LeydYbCVq0WWQGLTU/U268EtnW3QKlyGKAHhcgo90GKJVKdiskoU
2VXnrZ/uSejQGiboSVJRhi2XDZI1EoCTFbfmjgmrqnLPWDQxRwoo7S7hBIBi5kGZ
hJtH7GaKIm0dGyLXC94a+XUHjKlnpn2qDqQAOhTnvG+gYn/PEhaLBwXvZbldG5ZQ
zfeM/Qgisbno+no8iKWzTWItqWE1gRGs1P10a45KwfaM8M0Rtk2KZbu+IHQcItgC
zXeH2E8Bsts9LlIsh1DluVQ9YHJljy248DbwokZxJdb7H7aGtg0nBHisGezb3gMF
l9aAC8/c3dJAy5n7zfBuUTQq+OH/6NdraTNCVz5Vj2FLVJFfb55B/W7xJxzC5r3K
9S+4uHlSD/5oOY3gHpf2UQ495/baf3QWcV8USPuFXaTJgoLGYzj9344nEaaAPoar
F0stqfKu40ndrda/SfWZwJr1MpzDmPDphwqGbVKYkOQQFe3IYwX0aTbc/8cLNol+
1/7uCDbQRTkwCybpLSvspK97Lk6q6oyvLXSoj/Dr7WbxjJJl9P8poxDqqVZI/lLC
z7d38F0XZ1NojuC5yJwQpVrutwWzFirqkHdq6zyDM/HOUsrQ4667YduA6zF5DH7F
AHXvOe2pP4J5GfOQ/ALT3B9BJjBAjOrUFM/cKGgIMOnESBrO8jXRI+BWFUmd4vw1
Re2G3zeNE1BxuSecQiXCISk/fVMxBmxwgdVXZujy//lhvUvDMkNlftQe2UzLC+pK
QFoolvmMkieQRAhNxkzLFpV5+C1sAqpz2MSCl36ylFUhrMjJtebpU+mcOnsOtcyT
HxjND3V7KnnVPsryXUsByNCBWF6DEEl5NncyRpWFQazkpR3nDdb9VTRHD8gscfvP
Yi1s52rRkWPAkteaMnX81Cy6gbeNEy17/B+j2cUIpZFvcCaejdu/gl5Kl8CIO5GQ
LDaU2VWVQ3GYR0Wue/4aTQFuKs2VKpYGRGXALRQRxaIe57CXt20jtV1SpthlbPTO
5OVGljvxFRW3GjyMs3njSU30J3et2Wtw/aSTgjT00Ul25ZKHlhyBcHPu9KlQ3ozD
a5yuXoa2oCXWsCFkIkSL5hi2RkpbTOPiB83Z2o12fVv1r7+Td0iUbv5z6ePFtLj+
QxU8GZn6q7cOhKkXRipdR03cadzHVH2tuSyZW7BKkLHEMUE6IuHQDmY1OLGvIibZ
9TYwmJJDwkWO9aJujqHLTt05hIWMe1XOjxfbi6A3t7yTAfKebfSvcVF1DMOuvaD6
vGQCAJ7GUe7fpuijeSzQrHZx7569QomTw2sg3mzouSrW4GpJHiG69f87X6hCyv9k
AZGPrdF2I715x1AE4fZsq8FQZmGdQ9jcD+yjs4wXDAPP5avYisGi0AirqN6VHfMb
D4sI35smi1STwUKC8qPwmdIPj11BOQZEU8Cc8A8xGku5eFwjYqTHnc8AgqZmL/07
oB/fnbt76dnB6mgc6aExhbLb2B1Y2I+JRQqTfbxJY8WchYqVBkLYf4cooxR3den1
BdifAOiM+Tn4g/s3QvB12IqkVLFpFj+qwwvwQ5qpUqa3nCy2OH4gakrGIvgwXM4D
l2jQAC4Ue4m94Lpvi/w43dxYktFAs16pqr6JlnJS7LJ5ZShLJEsGg9oKGeaYk2lq
u0rrakAfJxWFqcxsJ+EmvYJiBGDb/FMix8LADi+0JTPGxoohnCPUnUyZW8wqUXnZ
QmWeT9yk8fCVsTvC6v4UX+rpIesuK2fbQo2PWDo6HPnGgUZ+cmEOyJw+dBnHqLw7
nsJSxndm5g5mQa0iSWavwhZtyZ66RC7nvRFRJ032NLzpHZmF9TjRMngeipvtiHdm
BAvqB1hHu+t8sGvgHtA4hWdEFKZUf7DiQeLpZZOVsb2SuFr2rp3dR0VD/bKQjsed
aa96jMml9MF91ZTmYGIgojPteTTiQCT6l6WB5HC/c+nuvBc4kEaZQFl93u2Y/nqZ
iuL9syOX7aqkqbGRBOI1pVv+faZpuSzvCe77RI1KROlUlVXB7p3Tmd39uvmHyncT
+2JVaps7y6550dDtzgrU5kReXioiZuuI0NVWkneNRvNq0mfN4nz6JnrB7JtZCvZj
SKI5nH3gC3kPf7vtVqzQ0iDNMc0TA0hym4XdvPL6Mhgtu0INwtlNCUsyiTSQs2Q8
kbTQqCQyjq7FILLD8v63RfylhNtuIx5SBWF+diBbexeWEhQ+rThnXKY3YItCMFG1
H8h+e05pBad7pgPNMfK0u01WeyVvCR3kQrScQlwDCQno2Oi3i23VfdLz0djHBmP5
3YlX7uZADkQccVIpkoWM8ORPzYciqK4/kctkuusTsSzDF75sgdwnrbyseYbARewN
QxLJay4kT7R6FCfcUSNmZvmEOLT6NxctO0Jc/YPEgzVQJ1LenHpPfCBxtB+PKF47
CE3m0PwLRXuac1+cwRBUjCEw72UjsDIA0zc4H7OlImjYL+JaJV+U2CUMOptsJPhh
hTClQmu4IFuPjDUckf2wTpTpG797DXmdkO5N9jKyDn4ImKeZj7czNY1QUrWCBapp
BOXv/KLawp77X8HJcDKzHsEeWzGV975QEio9Dznnm4Bxbp9sNhyLt71FPJFNFrLd
GOPErRSH/yugFCI3nPB2qxmDe8fPFP2ECFt1/pkv0w2pcY34TA3BuG9t0qvTKg/Z
WZ7QW/rCqrHZjxBL+LtpsejCnbd30yoYfTNXFq6UN5BiKGqbHGFFvaDhLYNMaJwA
9HiQZ3+Jsvyn/nTUu8o7vnMl3Dn/3MBZe0mm3ky0cBrNasinVve4+tGrEK3MbXtU
a3E56mfInAXWGG168qSHVfKWjXWsNLENiXokrmY9Th+9Yv8m98iRSI1O5YKAtOpU
NKiFhBd0Yk03R8ROUl1r3skLy81wZDmIx3GHlu+vLnKc+Y3fLaecVOVu9nXgK+bp
sB+EsUz1jM3vG2c9vXeJN/LVer7zqUmsG40nu6IpFYUTsQB/sCxPEIjLCRZsBdW7
PMqaZD8GpUhbHweyfMqEPn9usozOtHaYPdqsVgRg643BqC1CgXT+cdGU5Zcfttsj
8EGpVwGWIb1NWcrQJzIbm0Wr5XwxuYSEVe0AD8CwCcOxBE6wNFW1uCnuQoNjb9Sv
QqnDXVW9o0MtOSisUkqtZnPaavXpMhmcOADDaW23pvybruCimKC2RzAusv+smfbe
EWVa6oziEZx2weBSmqZp3vlegZNb2ttt9r/2+imd/csENOKSBabRYaGwy6iqZsVI
5//sO7L3JtI59YQWsat2jlUHh8z3MsAYiFwivOE0+U7+x7pot9YshxOiN7/O/atd
KQP95dmgn0ooIY3k50KEkGhyciK5hxjcKcblY9KImv6vc6Pey01YBetmlMcR4q9Z
0HhwqVxQbyY12vEwsBBSRYzarg6tLZcz0vGNk+4NT8W0UU12Z1iMAR771Qy1Vydp
O/uoEisQD2fV0/3xSoETPTQp7O//C87+Xf+6vewIxulGy/Ah6h8Na+jJmY1BjnpX
xbQhoqoxoHYcqwRCEyyvAPBLwuR6RUNrCNrjnKbC3pCu4QXgbwrUCtJ2E4QvqOA2
ycDa8u34ctqUujLq72q2UC29bRD2ED26iISSekGUmly6vwK5HFaU0c73IPsw0MoC
HyVa/eS3/Wl9NSxfVgQgrPkcpP3uLPFr6NfsA9rIY+/Xmz3ZOs8nSsXvr4AQTMpB
LPG5IbyTiIjlPq6xwwY2+j2yS2VBGximn9jBOmoZmLFy3OqetrHc+3m0Q9rO3nvW
gU7z84KIvtUT3LliakH9a5BIEK3vGbXfxP3z9Io4iWqWB1hY98blPynbou6wOaRt
Dp7krordjS5N4gwlNfF82G7uYxDXl6Uv8UxtYxdudOzKTyLNr61wED3zezn8pwQL
geR3R/Cc9T8+WIYOyXY095v13I5z5P4oIiNIc5nikSXAgeGHuovxoe79xdKMHHKu
6x97xW6mj8F7buMO1ypMGTTKW7EdsjvS40SWaIgqzsq7Q6Izf3vfJFQJClyk2UJn
uHWCJkabEYMfqNdbHy/nvJN5GJJ2mQ0X41wuna9H0mn7uPZBqpbw5R8FhQnWskVl
Z70iSJ151ZiVytDPMW5h9koOAXShpEHX+cW6plSNsn1R/J8CTHnajERRPbbAzlQF
sZEOZI6e8Z49fMNdoQzWW8pPlagTCHLGIuLSrzpblJO4dyC7AQfbinlhay+gZ0GC
cOyuYLOG1RU4N/w+HQIsLRJY4KnzlNYnfOvGd6F3u5iuIO8jCk0dyOUqCwpy5D7G
uKLMx5ZeorDZKRxIkkkeVgkbDzuVM4oRVHCsN/4hIYwF1R624oSoAyHiNuZ+EnXF
XQ3EVHUudau3cjlRIZmm6N064cb4Rj3BUf3Ngul1bawaU9K8xs9nrb1KjdO3MRkN
BkI0JcVbOrTWJu5UGF9XJ0VJ1dzIwiTmnDqflvE2S6MVAsM+Pu7BXruMzY68kthr
f3o0/q4PAuJy5/UfdRdtsA1iyRbLjsIvs7dyjDN7+CTSCKAxD29D1gFg0BI4ynQ6
1j9vR5gJFjxOzGjttghVWzXpoM0kgbtf9th0pcXRmAC+DshgRXSowz+Qwn/E54he
0mnqoGwO0fMJBW53wKiGZUQV4j4rB6pWlbdbuEKD5a7hO9LFrXZH+FYogtOlNoZw
z/Lmbae4qp38tqYw4Dq8mGWwnw7JX0HA8DkZNgG10LoPNg9KwQ1eYdKVB//5ZYdG
c5QAcBt4ag/B7jBUyb23ly8NUK+j7k85XUTcDt2Cxyr66x/6m8jy6mb/T72hr06N
/z4LOL5rE+hZeJPSq2kNkTllPOm5o41cXVsZcYdC6Pce2o6TZKKwoSFY/oy7NQjs
E7mahe9qcuglmYc4DuJSYVYy1u23ybJNtHMPZA3qG02POCfvEhiUrq5Ta28VXZ+T
em8pLaHVJMvgMlpCM9GPK3vhk15l3HjkFjVYidT9g8rl3Q0DtAKCl2RE9N/fYdBL
SVdf0B0EGXI05MgKqyd6luDYwiV2TfpA5dTFYTgUeU4Gcg6Wrbid2TyYrW249c5m
kNeFlBI3wSDmfCWFXaEtMerzJFO3rJsb8QN8C/92ItT7I2qRV5/af3JPZsC8bwXs
+SMpgisPWZ1oYMFCEotbE3hTn7TrT4cwp2VgQJq4ejIylkxgDzTmN6oDxZ2yBDRl
PjyxsTyPXs7bcVpch3c/m8rXzfACb4mv/2llT5pzQWAF9eRho7zZnwRD9himnY1z
Itn4NXBw7JnHN34pBrb6f7JiSKut6KnKkQ+/wC9znkvQ2EqvQtquEfAVl3v1Z+Ig
u5cleDvqN0JNIYD4GJ4E4vgbyGL2DZdcsFUFQmt7Rgh5WcenJzcqKEhBqpiVrpbr
Kjdz0Z6wq8YwN4ytX6XB9AHI3iforCZ5psIrZGq0TpRpdJ1Bft1k1mPPQQcDntnc
AHBesgM2vUwkq4PCy2Q3JStys+fMPgZYTp6Y7tvKjT/EpKWiQbH0oowigk70NCQD
5Eg3Lq0rF6E7VO6K6lwhY0bIBixFUQl7b1a4ag9NZ2MQej88pYCva4iAnA7HBpu5
c44+asaxtfbjh59/JPYewSGZsJwMB5uJC+ohrG6Cz2WF8oOcomVR7MF4Uin0qp/i
YOUtZm1GJUD87RjdL0J7XyQ8pxJDGRWrr18hsaQQoAMBE+Ll6YOqHSzls8euVP9c
DmASGTDRxY+uNQ5dp3XK0Gi7l1gNv/YwEk6W5punwncl2jclEM0Q7bMmuLkwESWD
kIq9QyjeXPrLqmcGTa2XjPArySqcfsg3NtPT7sxAv731WKbCZ7HZl7TIBLQzr7Kk
L8tKzRKiSLPxnIL6MD7U8/m4VqfS18hFJIEbQDezfZjCr0wyVP1HQAKHfc8SpCxo
wfcFoamE7+Nkej7MWBiHkIPlMTX2YHYtH0yevOzS+1aTIzr30sS/LEihwlHUuuxK
gl8xFUq+OH5QUkcV++Ca2VrlH2iN/7npJibkH66AGanrMyNVnWQ3JE8RO/G6us5F
HXE8yrDshFiWrFDWnxoloUNSlWgn0DPE+yskB62YJOUPp5JSsDixH0umrd09uCQ+
DxaRgf6SUv5VTSeKLg18NAKoQeUjhHJc7ydvAecLA1BxRpUWeSW1D6yzcWFW8gWj
30JpUP474Vlj5s1dWjH02CI85wejwlpz7xTa1h5fodhJnopIXMsFo1cFfBoCVNYA
BuJjAdIsD40x4dGW/kPT4vFTg3GuElmiWo8l1EQ8IA4hpTd+0+pvXTLE9lPLOl69
wy6CsUgVwJq00iUW3SOOsUd7E4T1/puT81CcDoqBT+b46cBgAqrFAFDUxr6wDAc7
UnTI3RuObPGPSzVpblp/q0ulB4ESOPUr4IWrIKBqXD8tcz6iX0w3Zzh/o8cJ1mRE
IuNfzkkK+oUZVLi3pvGQv4dXz3sgrM9KV2fOml80FZiU2mdSQP1GUbCN210QnT37
c+sDTfwlYyDuf/kdwZiqPDbZ/l0MRwCBQX7yk76wIh6hHOnnp4DBwhMR8cwHQWDV
1C11FLDAs0wasdt7VJm7J2fjal2ff9PRbEWks7L/BfORACQr0H8a+shNU/ehtFlZ
9HgWFm4tFcubc5amvBuGrsRBXD6X4kFj9o/cRK2I4phAh4G2dAu9mOLufipc1Y9J
RscKmqsB5RXUTvbf8CaMLSTCBm0+t/A32sG0DJ0N5CKUQe2ouyT1+gqQsu55pJQ+
LIQ21gHwSMzcbm8cn7akrZ72dRJuL4TLPUuhARWoAmgmjw/25SPvSGVTGE9S3Byj
uoB+SmXyN6EY/KIoEhxyoCNxPpqDIpQzYS4vZ80IwBL2isUyEnmowpGSO6jBybON
5jeEGa9moj4HrgXpN7CeAVQBxu0u879mgzzPOuoiM+YqiwdR8yIxeAvxZ9WM4HUa
OqkkTyd/HFrnmE3bmA3iNbMpac02Pj5vPzt0w618zammOfsvu1UBGCDLbLUZ0BNI
LoigRc8OwAYRrl6bC3PJRQpu+t0pxr9/JoEQ7gpxydmnFiqZXr8IsYOKx5Lxcu/Y
FGrbXwyCsnRuP+xdEX0U6ET30pnB6dokhJQnYA61wlM6YH74YQMqJbdXVxA51EP/
+/1qBSsIMgM9gNVBzLUT86oGD+JJAA4i7MDIb8H56viB2Exx03m6eyUgJQffx6Gc
9vnIykb1SDVP0cfvr9+u3zaX4vXShP34hGLKs1lcmoA30igtPC8Kk6icggp7p4SI
RnxQXwBq86EZOa9DAwP59wchPhQXXUsWqNZucJCZXwSOo1qG4V5GpFVzcmQ5w0mW
vMv6CTHyKIsR3bvfS6ztRhaMZaSS5WghEdUYsMN6xAPua+nOwtqxdBnEna8mLvQr
+haeEWPErfOElUBhS0xHLFV7UIo5GmIY0wv4sCvD6WYbOWHp3dFS15qU0Ai6f7oW
WFXbR/GW6s8c7xJGqv7ob9AOwdeocZer/GSV/fWFVivGaprrtAdmeHTPXF7gHKMR
9ojPRE0/lhyCnJgucUEDHUQlZSycFqaW0fgOB2eetm5ywi/Cr80ctk31lpV+0he4
1Bu2M5fySERhhs9XQx+y+FAhuPjEzfM1guM7VUsHFaideuFXvLdiUux6azgYkQjP
67yFvzM5Z22xshyEu0EUSAME1kmAxLcYNtfqVnUCaYCvFXHQDG6m+UxZi6C3mamC
TmapZB3dRfgi5DpAIhW45d8iozFUmNMp/fl3vphbNOZ5N027tB6z/XU3mibJIxYA
hf64tQZ0UMxLXKkwBEXUicL6FUnZiRxoAfXYj3niMapLeDjYdnbeLsO1gintTU4N
amhCQXfEVS9k1ZRhL7WCcxQyHINFB1fBznF1UOjcuEYUEp9jwkpo8GSEdXuO/lAC
nyhTp5gwe1XeAyMHWvyDsi5XSGZcvOMvmc+qfP+nJQy8wU8VlO3mMjYxySxaeCE6
T7kdYg7Bp/87wMzuZBMoOVvaX7geHLN34i4gSSYDeUJ7+UOHVq9JmsSp9uImCfO/
dWDfERCg1Zvym95hne5Bd3z39FSml8EfpGxY/omcC3eNbSAGdsvJo5ZP5A30zQ1l
HeLRlMupfYwHUkYBZZbWPEX4GJ4qjIl9fqpV2BybvCeAA72nTSfnO2OYtDVfRank
koWwjFlfeXvlo0MIx2Ccb2Wp2vreQ4vSoUP6ERfqBqInOEbwzuyIT4uJYLJrNYm2
PUzctYcAs7syFr64/eKT8onv9hwzzbMAZEKcz5oG/G3aPQTKfP8VIh10LVAuLTtV
8x+PCscv7xbCGCBkZ8S9DtphoekLUl4WOqjqdURgwKZl0yBJFkfG2Av3RXgn01U1
9QTQqtOgtW4uL0yNTHUeh9Svxet7YIPRH6MHh1JVFEo7NmpZZ4ZLAqkwqPFhknqH
MJ/ulhVVssDOyF3lJzZTOKTyF1lT4gu+i4zIDEO2xpi8eU3Qi12AsmemPzJ14xPF
N/7O9zoi/O/DFlhUd8djjnq/a+ZwsFHMpv9b2j147/NT5wTxZIAfuRbwKaapG9kc
VM3vrd8U+cCjavA0yFR+rOI/HyQ9+03Rbm+vrYeBrMS/GewvrXyb0i9Jgll09RBM
h44GlVVdufhROO2wDkyrORKLcR6QUYi1DGfwH2vac9bAz5SlXbKYp1lAFAkKIloJ
f/phKF+YrxFPGge7XtxqHSr+tgO1UkWCB7QbS6aBO5ErbuGv679GkHlcGowlE9zf
nv3TUrG/9Tl7AOdcdU2Pq+LKogdoRABz9lfd2p+Ur/xnVnfz9YVpK0vXbqnWfey/
mQi0Df0J+u4OEntxK5UhGCgUE44082DI9+nB3jJKK3NaVErFd2us5fiKZq+IF9oB
PtNk7NIKrSotK+vmA44V58dQVBv61moBvRc8hHhRRpdZYgV3O5PiTBkhQBIb+d7Y
sbbszuGsGwUjNJPSMXbM84qJyXKE0mb277z1dNaOXEYK5TyBYjFmjluLwqKFvAOi
w3OfGTy2ilmK3rkziDtDoFcf7/ok05t6xuCTo/xzPmomdAPMMfWPnykYkT9O5ElJ
zgOnkVGCacohSq8Kk9EzkaeD9fEKONW+VDJrgDjurHOHJUD1iuv1WySrgu7+gi82
mW1qVZilT3stFHYiWW8p/lTNyaC4vbJvek5ITQ3zRNqz8MaCAN96B8jw6Vm8bzyL
jfjZ3hiiJalEfJg0+lQ6NyMAy/T5eoG3ksk+SKduWGDBWZd5jZQ1czBiAsYZzciY
JoPR+mnimyrJtKyv3M8LwdI8EfV6uhQnx7Mu9vRoA2Yz1wQgRcV/L8QI478k8Ilx
D1rzP0s+pHGgJj4EmcaZwBsZDAESNs22J7/NLx2ZtW6C8pW6jCKvF8mS/B+7WBUx
vBjJCQAXTw9Oj/B3Bt/WepyFRGGklp31hT0iw5LvrgXOBRW/9iTK1V/+0KJNFpoN
N1nzcK/sTpCgab2PqyCdQ9sk1zo5XdGAbtQ2aHElM24a0ZHlB06egnDW67oEPTLm
NLLG9YI4xcmsNcdPmfCXE9JHbWrWqgjCUy5nZ2Leh0tKT6uR22rWiBWbQqMMPWQA
xggqGbXQ+80jczD7ABfmZJolIBvW2VxjcHKV/tflDRWYfOh3v5g4EcLSNVdgWhxa
bHPQJLrcJkGIbjAzB1u/E2wrbnxmmvyVbhNpmluoXDoVNz/91vqAYKN1WTkXVT/Q
PKRpAWgapnmEz1wH9YKPxKeexkzMAuqs/VEjFSewFkEiRPN+V0q7D9mXb16CfHKy
DQgwB0ihhkqCa0nKHFSEwkM+KswlABxVhDtoog9ck/T8ZXPSt+Qt9KWw4CRbx8NK
IgZWMEZmKD2qRaBkt/Rd1djRbBB7CQJluu1fbpGaxdKk69CP6JMCCCurGmhCT3T+
HD0nlODCrvk8ahdq+LM9uHl0B+BJI0PG6q+bWsKzq/Si/CBdunY1Gs/AUvAyyJHT
SFNEe2rTns9B5YhuNX5EOuqu+V71sJY+jj/hF468HgezjyTaAMp8rqEED/0hHUKx
Z9nD/bJ3EvTffg2IduBI6abnrViNE2l9QeVQfbUmh7hjLDRSpzItHxFDebZsXHkK
Qgb6AYL80ARkmEF2odPvND4B1pAOJxctVLhLXx3ix42jzeO+O+xZARhr2eETjggO
bbWUXwEoV2EDJyq9296br1JlGtXjWMVSyxN1qfyaueAqGU8dY4173gr5gAU0tzM/
8Zn0bc8WkLjfLoXT1oIIUDFNM2b+nM4p0YfFcAgx/wZgyCxpQ5RNB5P84TEmcIJR
DJD+9PHuyRo99z0an4O+pt2a0V59A/UBFT6VpbPGFx3ArUaCpc3CGpB4+35B+/m7
29uWGT7iSenXIAfcehog8uGi+9XklQyGmu8NQrj7MeA/orRetsIodNxwX+UsEwjy
AMwtmS+yx5kkJ/ReTQIqy7Rerkagh2jjy8nATHDeFWKEHOlMwFEl+vgiecv4Jmk1
L5spbyiofBUb8AHia25iDnpu7VwDRef8mMi1f+T/sI/vsckf6p95dYEQjjyJ50d2
U3z/hsN52Hk61Wz752fOPJdhigkLx78cYU8n8lyW1U1vEYXiKP6jYLpnjJW9Lzhn
eHSgaaHNeK7NgcdHFnWEUQE2tZOENhOY/06Lhf4srAeFt8w7lxckE75QK1GplTXa
b11bwznpbE3Zx9Nwr+XNg1+VbPuwLKM6GgQdMBWtGS4DuGgI0gCgRihc5OoMtn8G
KjTXQGxcJUBVmswEc0aPd1MWE11XPNnEceoNzZkmq0EhLqu29pwD82pRGo1jiN8h
DHqQWF5V+cCAxj42Yfss+IJfXCcwStOp9aLIDHFMHZY36arByR4A/m6GRX1ynzqy
JwUy3FfQGczJf6suqFKlcoelCBYZAWKhg1HPxf8HgpwMM+wZ8ocBwQjX/TutBFAG
pFX1QRzojSj9oXWDtoPjewt6d/RgBLp9g258xAsRycrjzls4mJNFvT8zI4i87kaF
rVXRG3Fe8CtZ0hb8QIhcNB0gPmOsvVpyYmRR7EXVI+kTZzKvX5ko22SR51LSSUgu
iADSISsoaoEMPfKosIAuUyngix/NQt/RNyzhPFi0GaWH16Ns1pGjgmGlAJT8faE3
orHcqWSFznEe5PqFhmXBtJJVf509M4OG3cFy4S9GjgFSTQlwJx2Rlv+ucBWOjAiZ
paOD9XcJIpnNwdBBr9LTCrM8NPHZbkgcmvQofLApD/dTmqnZ2DWTM7OpjIFF4WU0
lIokZEUeDLsnjIDbpQZBDVE0VBDaIwBwYSGCZD9CnyFuqssjPuu8lo1f6zoCw5ry
6dxOXa84wFI7H6AwJzJWTxO66ZRDQ2hRybKkYNIVUgBkfkDJYxefuycSYx5FYaKo
k3mHrXS2Dhrcdv9LqqEW9HCj+BiVM7ysvHGaEHpdtIqBssJ7kO6fxiJlp3ijwqd7
6lwQEQtI+7/18dzRsvJ5z/uolv2g6zLuo1Gsi9XglmNzEInMsjrM+7RXfNop7Vxl
x0gJq1LtokssxPFhKvY6SV60briTHqmT0wjNvXIHsDPZT6ClYg1+fPvPRxEjvMLB
dJCGTjHBL4UEAkqZ1RcgeHt+RNkPYgGxxsor8Yw0p0vyQus1DwlTmBNT5ceBpQdB
AegVMMbzxOFxZjJCC8pC7LLhEkkcIvHdsSgx5qokXKsyTocz4J80wyct2UcG5fRi
aFd9r68hrRKQRNPQZTR+mBvH5s+pfNplyEH5Fcg85H/3kyXXI4Ut673X6ndhTC6X
u9zYxpMkL40S/l+e4We6BTPVrc7j+PVczdb01aM2AJ8eBgp7gNEDzyxzKALBr6XY
UZe/V2fWSWcKb9QDyJwstj4Fux4CXKUanGhXKo0YqgrMo2BhvzzgKPGc9FouP5EZ
GTtS9+ZOCxyAjjP0K2qvHKLFRmp7D7+89s9gsE42O+zQWVbrM/aPwItkxwOV+FCM
Y+7s4KIXKTZzv5Y0shADGwXm8AwjzwIakS0IDL0Kx72j5iq8cnm0KFsixDKg1oir
A+zlWwOt+ncwST10s9tDMFFTUp5Tny3tNcQ5pUiYXkhEXNFul30/usbfFwMqYWyL
ukF5XlVIADkHj5YLXI0A7EAXQTFwJCLb3vReiXfJK+pkZtt0JO4uti1bLvtLFQZR
r8jufe28lF6SDwJYFrZyIXzd+GGBggPtOKm7TZs+/a1cU83s7+SXEH3CFczfDtM9
NAlpe0zJBwQLo1tBII6bV1tSj7QFtU0Ly67COPqp9O6zlzMiONjkO+w3iGzTrt5F
hLuHuH+9ph00CWWXVze9PGK7Axv8Ocdni/BtsaT4DGX9WyPbuLHzqCFyjM90nRi/
Kg3jnEOVZYz4yRgEy3TkcqMPL6tPu/NtlC/yPLAqOITXGprYc18rr6GO+B1fAY6o
SxpZmduJLpWLkXN4NmdxbOAGwld+LWsgO3+J6xI0MwYcShMXK5p7AXTJtzE5LkUJ
M2QxOUlanTTqFq+rmgZldGUb1uvLixAUKwz3D6RV8KJBBhZJsZUBeSSTFhRarXXp
NszpV5jY08KzagjIJ3mHhI8gQftJBqwjpUhEZhWOqDiZKXOW+UDSHR8GwFDF62xT
/S44NCDBX7z54MslOtfGTiRfQUt9EeN2garNpciJrh4eOifplSM/nKFuHrle6CYf
P5ziecXJdubdARGbtk0mh7EbWMaAgWj3UzX3SnjgSxfyPAqNSqO0FdH5hxpcnP3e
81R3NBzY4+2CMU1JRJH6j93hWcmOtgQrMZMf+pmgWSFAitIK+3vqgOjNlWqhCUBH
iQqUQb9KcJqGNQL48dMj0LlTHz+7V06cG78zMZ14rAZfAVXKPrFTxQHWZg/X3nlS
pvSrw0fJBaYbJZUTE5f/f9bK55cwaCw50sdICvCrVgf1+RDJ46+YCD8D7Q5NeoSE
tSzGAejdvqVyzxe5pTMykPgq5Nv024eRxPHAX0Pkbb6JCPeNFIH4hMN286tgp3ll
04Y3ENIy3rNIUOm79YobeZUPAxBqiteHDYoVo5hiHKuB7K31tdj5coEvmwpIYtLc
jW1zyOZrvSi7C5t8Lwn+ZChHD/+iEhxWMGzfTwTNyI9UYyye6Sv+szB9+EsYHA+U
Xz5xR0nZv9j5Vr2vgWpAeT7UsEchtO1666nliLC12slbO9cB8eZ6/33HQTn1S3+k
6Yh2qk8NY4NMrMjBfsIHSISsQTli8VHgBNXs5uFTmnI4zWX40n+HFiCGLrxFeUrF
RBtJUs7+xXap3sfSja6W3k1JAJuiImfGPlcqDuyBZuk2Qx63UND5YNVxZMkqK51D
mxobz85xABHMe6KySlYWH0/WvRubr4bwsBDObwSb6l9LxEbHFvRRNplG4ILrMLJX
wWlT+ea+r69x8Z6AepSQ7hrtjxdsKWKIIfI3LcOwpXxzsRTMYhPtpbp4lNvPZr6r
ObKJ4Bu/pRKWvLwf6kOZ46pP5IKg/pyeGwvSShzHobT5RTiEiMqxPQYh/Pma7X9U
H40wgTYgNmHcWZv4SCGxhC2G0nBKnn5JrQ/CLQKF41NsCwnNKbIidFi+xXdONUVp
d0eAxCZCSmHqoBljZOKWO9kl7aY2A4oeCN9Y//xEMPApm6X37RFkTXOZyBRP8JzS
y9w1Ba6OzhjvoX1YygPKbRahHmodsMnG0ibWAXlwLqUpbTScbqUmhuf2yTfve1VE
T1rsgtfhFzBLGaQ+ta7jPzs538Z8NAGd2Ec81+zFi5+gzab2m0CagEwNbBWp0Q21
Lu0nUtCxnyCgH0enybvQIBac8kKd6nd7C64IBUeXzb+YBIUwCTadVA/YoorHaUOt
ewOrdxIvu1gBEkkCNMuFVXdKIU7rKZl0S9JMLna9JJmmQhf62lP2p5aQowVUbrzk
EQ6mDRovUlazuPzb2trPTDkDMJxxtYXQp45xd6oeX3V2M421u0gQc8E9pubngN8w
dIbdopUONNwk+IvP9J1K47Ntg6WUg4amzWq/UpKluvyguiPYlE5MgrUxUYGOlhLT
QCIjsIe1zi8JyQHssdJBeNlzkQcwTbYyXvKmSyb7J9TVRrd0U09d+pbyfGDdycvv
cr27e98hCiHbZmBgBS0R6jHpvAw+CyLFNqyoHe6W9ImJnQzvFo778A5nLMbfoEB/
zLL1N1+UAmTa2AhYmps5zyCd2l3DA4Sp024bLYj6ZmBkiQMRuNRJvWsLigQHZMm0
1RhNOhTW+s6YthBrNjiAwEqiLqViSC9s6NcpfYgoufkCVHocwb+EFyZtCbOjyK0k
ZN+QPfR5hAjyvjHYU6uciUopkBIwyVamM/VsWjNawSYOwpO7Zy2LZeQ5/H1cm8HY
ZPogW5DxJravT6YnlJ7BMgJW/CFjCPCkDB7cMe/GttR8tZDYhcjhmy9x0OVVXbUn
BmQU+H64NcOewT1wwMTrDlZUWN5M10BGnEmmb/jxnrqHw9STWx6opSB/cahRa0bH
1myz2eIGhuce+Z2sTnqpODwxPfEBkB9fCRONaJok8az+SEmznSOXEhalngg/dx7g
aNWyIuaNqgo59fVNBLqIovqgfZ4JPEyodpWU+njecVkrgkySJqYFueCZ9bI05P87
2rMZdF7T1KK38gcLMKBILsv24oy1Y2upumSOZPJkWD1VLp/PNZsoNJrJHqaav9Qk
fuupR/WfzzpCwO810eGYbFbAkvLm9PYtIAl4Nxz9DvcIoE/fQDn+spZIIBFyXY19
O7fwHk2y/hzHJg9IuegY/B/1L1Rfadv7UIsVduVXcfO/NU2+USecHD1FR0Q33/yE
17iDLYyIQjqxqBEJZxz7lVByoFdQhV3E2lvL+wowbiVe821RHpwhX8UJDWyLI1+5
r9+tvkvlPpaHX/gTHIIR5oNxHfcUDDnXiwhuDgCdDgqFQMhs8bN5Ac2C4uhI8TGo
TWKZu7U7Drwo6Piahv1+MK0FcFm3t1vXAlzVTA6+zJlkU6gTXiA8J7/v1/SkW1hw
qG5/6vDL2C81LP6QsaaTlYc2uJaVrVSjULilsI58R5tPiL/BBnpIGXZows/m5wdw
g42jVFmsF2vtwSdllv0dobZuhzs0r6+8tIbdSjUcamNsSDRtoY0jnRMpzsv7UkEF
iTMlwyfF4c4Suvg78OcfFRLSMpzsH4PF7tDHrixs/qvbG6O/93/WetLFOTWmqOBH
AhJWcsxo3cebzo2sN+ekgLkuhTHhZIFrxSMQs0fVOrBUq/mUkbTZHAx1inQAmErd
HKqluyS/yp9vGzkALW7N/uVGC4e7RBApcLSJUCo6obAkMAeJBFPIDf8z3VYmm5/9
GL0/LyRHVE7tWHw4FiVOpsIYgW7j1D1gFhLkRdvPzPg+e9yVyeMpI75X7Ejcdj3E
RCoBx/fQ/4LUgOvtCiBj5e3b2Itqcvg+M9w5tuIWUyQXaXeJ/jquCCf7WjkeoEj5
XTY0YTtR5Ve+U16tAWt+ikPq7vvIdrxQIf0zeGAejSTXrAflZdb17W5yfPlqsgSJ
tsqnvwdXPa3as/vymPaSk8zKtNUC3yGPlV4Vrdhw8hw6XEKbOGO8rnLg64dm7OOT
YN7XfmjIUdqC4lKMQVmR/k/p/l/1oIy2Eo3pF2e9EBSYjA+o0OcTSgYGfuATRA21
b+gGcGn2YUls+TsiVAh6Pav1JGpbkAGsnxcOtjhIH77chFU78GsmT0/yuBqL2meS
zlJhmK2RdM+1mDCqW0L/CNDYGeaOb4BifOYlmx3RDw45r4bdrINcfrryXbcJy9Qz
BKgETqICYsx790iz3rkcgQdoFCmB3o2MFo+u/xXkX6rK8BnQ7n2KT6iglAN/ULr+
V4KhMO27hqjIi6qKrrlXiuvkB18sKvEcQ1LZY4qIdBEtkS1SoZ7Wz2hZHadaVlBO
murA4oIRC31cyptniYvn6VGYOKobqrEFoM1GlOT4GQ8qOuuxvvxCkpNRxXaVWVxY
Eb8Kw3S+tyu0OSoTCBVesc02ZBZutA/LfrOVixMrX8OTdfR2bgRtM1ZF4XLVBJAb
L/Sa87zBVp+ocmkHgrQOAcXtIJ0vBe6Uzh7x2pLzgddykXlWY6rvJpAQOuClzz4i
SwIVaOjWFlSkoGiSj5HxJ2Li1m5s2QsiPelKA1Las3NlNP1GoC+PQOA6s5+cIQSw
OEaYMmpuDSLiBJCUOkwmmm8F6ya7fxFc5i1DpXwuPzyttNvLF2G8GQu0YMAWboHm
6s47bg3V4tnUWZMynau9R5DZcrd/+NN21i3A8U3u6OMfT3m8FkP/ldVILHio9roO
jvMoMEvR3l3oU5A0Ccy/JEPokDNUtUi2O2KrHmTGNBo1z8QQ50a4AOb9DOf5mRMJ
FIOFjW/DmUbWpQvUIRV3re30uFaHNI2XbMC2w2BE0UqmCn/1e6EW/hq0YopfzZiQ
XOkKwieZJHLk0ZKiv9ps7IPrId9i+Ijk6n1C/I4vSwuspluU0CE3kSkhXYOkfEAs
NMpQFq6K3/MDKiVPp/9ZMjJ3r4/SoElkHHflgy63SrYY6E5GGMUcaTqqsFNg94vD
3963Sle9Oxj5yAK2qytE3ptQKcb3QMbAp1pZ9LdfnZw7LriOkSAi9DK2qV26RLVj
duX3TA+86yCVwzDzSjbPXrCNJqbASZ5fnI021xLaAXrZLZuFu+TdKSyZFNHJzWhp
M018ScGrMpkgzj0o/1P1rYsZIGnQtZxWGkfOdXClu7qAD7D7QpEGlHFHDahFhW/j
eDLBAkdleiu14tgRz/Aa/N0iHfUCQjLi3GHd+7H08xCNGMO34+ZlDBwqlrc4V1sp
q7U1OFaRYhMT2nh0CaGRCXoipRKcYMMAQpSJT+Mqu1BnyM+Xhndnmy9HFwA8Esck
pojcEQsJx67j74w20L7qeRpueLj0Yl3ZvNGu6x8FxfVDuCnTX2k4E941xclaUOdK
U/Wl+ZvRPO/GDvsupEyDbtby67G1eshMYWw7MSneuG+Nun/MXKYVlOgJsvgObF4D
M7eUncfKPxauEHxQiBF0MhNtwCZx8QV9LgBdoE53dGVTJ0ctFFfGK5zdg7mekhTC
uXt1FLLsJ1ermImit222HIuwn186gFow9XObFaUhSHrKyrMZ+xXAMdu9EUeml0ZV
Q5hDHI2CgKmrc2s/G2CXFyOS7Ww4ZC59F2IT21dfVL4HEsBcFB+4kjy5pbYW9maR
A9q65iKNZhaRslYL0aVr2cD07W9VjsuF+bSSp8RHzf6CoaKcvgzv9I9xYUjWxSjd
v7iZyn+7jfssGoaOOiSjEiOQtOfK08aKVwASPegfnZLfxPkHLDqmDBDDtdhn6ctq
KieR1D1Cnoyg0hyidu+VyveaGPjbqE8jFnG/8/BCXHWAqxjUJU4oCet+Ldp+Vu26
dpD2WLMcsmTs11J2Nf/WrxXtzARfaYXLz7NQK3I3SVaHwPAcOTEJU+5O1ECSKnQy
3sAhKzWU0EyOHNyDBjmaqUcBRM5stzWCIk3fQtm3Oxs8jnXecMK7/dT2qd2T0nKQ
7RQqXXp4AZZjHTec/qhFDXdkBN86XLo5+aLDu6abkSqvKiTvzikJm8rW9ThL9C4f
7FCx9/yCPVH9X33lgL+NNKgz9o9EimH9km+Za7t13IADvUGp0vUauy0jndCo6o7+
ibTFRuLtdhYpElJesc7UOV6FD3+dTQvPsZMOKOs9nTPvMHQEo35IpQYHr3qCp+tK
dXK3zZDKvwz8RDYBZK1wc4+DgABqo9ST8Qln22WH2aunWfcwuiaU12EhULlzV/De
U3Zi22/WIQcE80RZW32W7PaQYNXI7DUGhhGx9NPgPo8e6HVTRCdwaPuMm87rduka
EEk8sN4SvPXUNIOpQfbDaSRQSAPKVGmhuEQZW7CYF8P8uYUyB/kxEZ1PFjlff1uS
X2DNkF+Upki/o6kLuFf4g2Lonc9K88Ol3Ylq32WoGMjKCoWi69bJA4kng+kzq0Al
oYakwvn6alJPeyXnE3cD8vHo8nfZtfz7UNTdcps9BGlgBoN6fcWwKSU7gJhnxKIg
/j9aecXFImYvLnGV8ehPtN0Xm5K+NqeDekzxwrjlS/jY6Q39R5hyUD0qr6hYo0GU
cQiKyonkcoE8dR2OJ9uOPPGBJ++a5wUH0As0s0mNFR5iVzmLcR//gCZu36RskWoY
YFETc+qBX/0e9OTACLU1KAgZbFx2IEDV/a4PJKFcWirvE6Y4HqRKRnUFPpadGHUx
uN0AeoBWVCzGrNu75NjftTUE4i2R0D3IxYexjKJ3QJCkFuvXMv49o5nuTZibVq9R
1Sd2wS0mlKdEBUA3TdrWcC28KrJnEdHVtuhfonCJ5FVdtszOykfuUJFW7EBXDk1z
OGWuX/i1x2xBJucxe56i1UhQt8vDS0nh1zfqEe+sUGjCJzXYQnlGnhc+MuWhMnBC
sNzF0xlk4pJ2Y9hDx1DSoHtEBnuZrpCK3YIVxArMbnXKb26+wJxfJwh0o/tLFRNY
CNqeoxXLD4BsvBtlocJSHrEkpYPCYn3+8MQuCbe+8mTlba2n9q53R5nVHDxgsCL9
9kCsnQNLo7h/U0RCmDfudvjCia9gHlneVQLMkVqMVWyzlLf8fh4h5atk9jIDay72
UW0m0Hb52uj+u2nozlk+2hACzwt/Yfz9WR5HO9OKAFwvpLcBIsaCXJxKrbSMJbsj
+DFTC+S4gci1BzRCxCwDnTiQ2YxHzHSN0CL4e4dYru2eCEvcOtduhSIK9UFGBMzq
y2g5eTMlc1nvqPtA8f9Qu1kVjDUhmjejtBp//3YPyd0KlwCCKxArkKNfrd3TnSc0
iC3vpXqXhjk0Ltb3No4wAx5PmQZlC9g/rjyssK4LqWrNZzTr3spnQDAdjVvIxjkG
0y3Lu5S6g6aFulCBTGhBexo+roq2giouoVb9QSy54tLKnVofylD1IEZz3FLUIFNE
jDPxIjMdOHGmalchj0n7SXzLTW27Vrv2oJiwnVGamyRTmFuNjMbWHhRa6mOWEzt5
MHWG2jjrhxAvhuAZEDn8xqrcKCWvWNGHZipRlHPZtk19tSMI/8gHCDbONZNkgQB8
HTkk174Cx1N7etVOGGiHoSEL2Xxvc9s1fepgkWJQlr2zn1JogVG3SIBP6ueqvHaF
zF1fMTIQ37oV+S616wkGwDTQYst62MMsK2GRNyl/TJxQgmuGneFBYmf/sgjm67kw
Y7reKemOmWYiQcFcjtqr8rm/jm2stSZlMbQvPIt/nnnUbNDUfyuuqzrR6SrPitkv
waWbB8LE90jme4iK7tBidftIvLo8Ncu1fepTI7Lgu91XqzF4WmEo3WMoLKzIEDj2
0JDOZl434NGD7SZvl33UP7fzQtgO+XnL7Qk7vtg8SrcnE6cKbm0gJEFezfaKqskL
UbwS+u6JCDRCJJXiCGv42QKZhe/Mo+LUSr9lUp/eKVQ0Bzl13Y13aB9OS/EKs55K
vJXXUYDxvGIHSn2691otmo7pCkNh+pCnZhvuNMpObsw0JcI3c3lmj7FcJ4YFP5oT
8+h2ujzHuZGjLHFmnOwASwY9uaMN9jCjyBFJBizchxyLiFOu7UF0XG4W4mCnjQH5
xIyy8Twqactx5MoYSrKYdis5EQKZ7EdUAoJZfDunIeyRCFXNk8hR3ffKK6NAbpTi
+mJ1SbHthjNJ/4UVogptsWBeEqzPLTHtmDc7W391huxIlYs3SV1GHjf92uX7DVfh
KFiJuPJfFs/mIohg9S5sCSQRWNL8WJvK/gZMYAUEgi9GcYFRL8UxKf7cr7ZcQOf0
Y1lVPIuqLook6Z24ETDZRSYFaMinO75aZD7rpehubtpPjl2iwFRxOKRdkIgKXn0d
R85vogXsaYczrzEMX1Szp/y71XYnf4hL1kAICeULlqeNZfWjdifdziwRi6OmPK9k
Q3qVntUgcA4mlUB3i7RqsnaR3CnFi2ZBzp2j+HtM7xtoR2Dcl7GFbZs9VegDTRc+
MlYrVXwHgDk/M8vH9urgjZb8RJRsKUDSGisC934lCPQbADOhpRSZEOS1nyCSAhuR
8LTEcFE24BaPDjQuAo9N9reXLdDAtq6BgE8iiReG02NVxhhN8Qb+MWzjRJmlz57D
i2SmC1byXf29zWK4i6L1x1yrOYNNhPjTpgmxAo6beSY4RFajiytlE33rse8+yz12
zwk/ejkf4TskpV9/Q8erZxlQzNCBFdKjOlWU6r3ReXITWcLxJrOZZNLoJIkyUdg0
ekY/z/JXNaYZHM/E3OuMdTw+UXamqqwpR9bjCmyDd1xf4st3mNkjKTdVpRvqsP7M
61pV87euRt82GKiUg+DkHeRegwwnksZcaB4LDyFXu9yPaNFCZ4y5W9oXIRl8EA6r
DqATBfOekkYuQlwrx9YafFHH4IvyKTEc/zYpFqL45vmWXsY5rmosxgagrfhV7aaV
wTZ/XEZsrOEvenldq5C+SHSUVzPMXm0BV+3yd6FPWJtUMr/aS8viGyTLjsgshQbC
9XXYDEAioU3sTWS40cecfcl+jqVIGnmE7+2298yuHHrsZSKOAI44QwQpshXTH84N
9EIJZ7UaI1D9QJg45r+SudBE5EgwpKxh5dyT0rEE0Jitk+Z+VHYP2JS8oLfOoE+m
CzJOY4YP+iKKu5CgvfLo9hRX6sHAIa9jNWrsLxRy2xQp1wH8Via2v3ODm9zaUTaQ
8aQ2CPTGh9Nj5BrpFWJPxLEmNF3TBS2JDvkU8O43UJOgx59IeHhTiz9eCJsTer0Y
lc/L8zJkqeA2vfjwG6VONNt0E+MacQeo14D6c+DZW/PT9/Wx3irA+8AjoFFtCX/4
/r9N2BkA6ziUKWRrfs50O0Hm3MfsTCImbS1wRZJB/mFFtdwgTTlGKkwtBuEnmcEc
hMAbE0hAR0br+mKwDXEzQROiJJVgq9r/Rd37qBgD+jg7IMGopmaBT3f+DaIMh6eT
/9SROVV3qPo9CSPMQEa52eh1MTznREY3OMB80c4lPXVKMwQMmXkqQ/UBHTOYpJj7
jILRLf1VGbGlKKVoo+OqEXd+/kftYx2pcp7qI8FvNMg9E6H6Nzok3mu9asUZxyLn
3TJ5OON1CrViUUkkWXU8gNzcW/hYjszDDWcuK0nkR5hX6v5GsMioChBqi52DhPTU
jFWt1ccsN0n3IpUmbtulWU91eCnju0k0wvhIPMK2t4E8Y5K29a9IEICKIg3UVp5F
OmOvYmmOCOAC/zJexxnATZKpr//vamQyZV8ER7OAPGLRzjxh7Q/whqvJZeQY2b8z
fqn9cOCY5pLMpZ5Qm9f+1GPxJIxHrJHIuijNIJKxcLtnLX88Ow/aQTVk6S0QXI4/
z5hfmxszp7YtIoH/mXlAqsXFyKXB8tVboXea5jk+0Z3fIlmqBwmXArQ6l/1dZF4R
O2gYQezukTDTDvi+FwHhjmr4uQlVrxbQfDqLu/Qlnzsv9CxKyt8esn1WlsNlxSJF
jQ2DBppyTbNWM8RbuokRwzrLxuQQkfIKjuO6S2nuZ0NFeZPzZQo2rww9H4fE0c3q
FXUVjj/qF211kPb/v/DiqZuipoQAHvB6uDg5yXKLSJk3L05xeKKnSrcmiBpEOjWa
R0MXkNqWoo2l85Sfe4eK08ahKZSBQPaSVN46VvSkzjzfoyD4tm4ST53aEdzJ+MH4
+ZAOqsa2XbEC7HDWtgySgEcRwR0PGnBQMbWhGWL7FWCJcPmxsq7YfDZLtk6OC9jc
sPHw+UkwiCeQTMIeNLgDenhUGUZbvNV13elHB6cAgPhVTRshbXd5ZqeBqxGUzMbT
FXgsu8QbIXmtEP4vrctNYafprna5TqJxvxrs632NwTDvIxm3gE3IBilw26D8miCa
5fxDFI3APic87Uk+e6OuJTuS0o1VMejYbu2PGAXYyWYMOxIXXxk4a9lbOgswRwz6
FFY4/6mnVzK/xGC6nacRKBNfHy6Nvz+QlDayMxhxN814oKxCY+KWG24u/RoiKnOf
J+PeqJig8IDlaaF1/DrrUUiFPOSDH6eiKz4lQLVT6Ub3fij9BjrGDsQ7RwOPz6p4
S7tb9bqiUPL2aOyLP4doxVPplEoueppuKLnlCs8IduPczvH9TGZKKk218FWxgbim
0/9evyDAqDvD9EfPJAUGgxFdXUHQNBzWZtorY0zJUHpmnAW+Gw06VnbEVWCqlc+6
9GZccwiq6/ZN6npdpePwbLk4sTf5h7JTY5oY8VjoBWzOHCTo9DaP00rgqUq0L2Ko
U6dSHdI+Vl9WWJduP0x/lZgL95zl1UhsV/l9Jr6rq08XHj4og2b6RbmxziaXapTk
MowSAiJp7T+TW7pH0xpGX4xHOspq7BWPCtqXql5wlKs21xcE8AToROsHLmkQynUO
OfhPzjhC0KGMZc8z1sxMpHuiNg/MKKZN5qg4aEtsuDTg1//bpizycSUumCCYQQsp
NAonQ4VoMiBaLGYwATPHLBEz0hH/ayETmHNbah87GAqB6xSQShb5xEqs8M0p8oKi
EvbRt+ytaWScFl4XQqZgsX6tkcsMzgVaKvpjnoUe2jZWtqSSKWoF8OZxH0jGxcPE
LvWJmaS0AXgklA8q7dn7IusKEWbUJviWksBSLwP0gn0ucJwqyXmQe6UMPMfsDPHG
+efoYBqv+LP+ulcz9XWFC8zqbknhu7pd8VmeC+GxZf8zeUxqxA5QxP+G88Y57Fmp
n26G1y9DsG6rA58u1PG7K3a4HKSlDt2mg9ProXbR5/J5MVoL2kWo2TKI0/Lr9Usk
/153frKk2xsxx9EXFb9rJpZhV91IKjI/FSrh7x0SVdvxshWXgU8B+J9TmNyYM7XQ
AE8wsInRhEkgEE5z4zt0OQCdvfT1sdw6XgccYzYO/mrv6UlNwDbek1Ms7uwiFOwt
qRePM9wQp5xoj1lymUJ2/v8YcB/lVh6C/Had2kdcfjcWHNEXHBt+VgnFEdO68NGC
nYv5nWgepffq5Uz0PQU7lA4NaVPKs/5uawQLTQu5549O+MO5b6XpbPIq073/iIdr
I7B6QLzSU0P3iRMsoeP3EP6f2/pxRjtOUSFHqBO21/QyiHtiFHuVpIDr+lNWOXIm
jvTYJVSDz5E4P8PgRfy1PSMJwO1gHwsbTdjGGle01HMrhWzJNnzrf9rI1BANGDCA
3fPRxPB1bQ8I7c8DFV+EYZx2a0b9Npu6D9Bfi250fNCmM/yF7qzWIsgwI4eHuIB3
6ePKNQMVx7Nxr/7u8JwJOETaauD91BHSh/U47clLUMWqFxwP2IQAHDVCN0vDR0dm
Uyq49c0EqOBVEMUIs/vmZsQUJlMUYzk+QSmDEIw80O+teTvqqoX4udKmuE794HEj
Igxbjo2caGV9DshgpdRwB+nMFdsyFQRXNpWijTpaiZZiHMxi/wNVGOjfwE37auwH
J4lAFmPhELyppRgjA/w3OrPba8Jp/tD6qwsicJH3yA4KOnijPz+OhqtZS0ZflS8K
UlxKPkZdOad4YnEoKJQf2xttxunbaKnPsXDebU9Bb8ZL01X2L4f3Tj/pkQQmEJHJ
6EhXfWUCjqTdYoBB4/pM4mGCR/ebbf2n6AzfUXgfDnrYjM7I4RGqBEJ34EXAXAxw
92J/cQ1lKv/GImtyV+/YvSfXl5XZ9+JhpP2N/7quoK1xdBTR1naaczMgWugOcEmI
Mo1VsA/RSY9zZwI2Jqc1KVK4GyDfEupSEtzqKpi9mdso5kf5a1cke3kI/eBk7DSD
ZFbmYi16Ds2ksASQwKwyOE0PGgCWx2YAtRs96Jn6acQjdwi7+I7ggzbGujnmTasO
2RslsOcMeRy0PDpAhGDiDMhZIEDJRpOlVp6JCFC8ooEGBQPjDfGejNJy6Yd/NwJ1
aF0Mcp3OwYB+/OgJ+7MGhaF/ZAyAYMUIGh0kWWu+D/jGtMe9RSXxsJ4gsAmFEa20
GAx8TACU1FQ+SpfAiYS57UoBs7tISA0VfVwrAFoTIPr43XLxPBO2JVisnbx0tqWG
GlSpYVgopyd0EHbgRO0xcrDbvSjCFM0ih7YGDjf5KpzRblnfTDsLRu8q+mRNSazd
EB+A9ZJAR3KW/ketizfCMHbE5a0q7n+xK7BbyvNHJzGqZzhO3uLTGIm1F6zFv5rc
aNO27wJOFFe6Jr+Ml1AhLf0HahlTJwQQ/KUHHijXGtuYxyeVhqNEMZR03zzsxIVN
PD6wtAsvI746fPJd7Bn3FQ4jbt+UgBXGqD1s7K8Eha+AL6P0xT2/6BEvMfxv+ehm
IZ86ssjnLoTg+ELj0jZgrQOieM566xnM6fcJmMUYX/SRqifKWZbQRSEw5bTOZs8U
WstaOGrv4UogSa8GbNDBUk0l5iiHdJUXDlNRW73yNDFrNSvJ9rm2Ar5VzaexkNIq
Sz4lJLo9GNwO0NaKQPnNNVJ+NC+hyCChsWHYFn/J3mM7hRZiiuCh8nIJqvkszoFb
I1nZ02sE+cme3yyYLbQ0wbX9pK/PgoEiWcO62vXq9m5lYuaA0SfCk5ceQSrWN9cU
mL6iPf/kOPv5mfEEkdldRI6AmnOTGvuid+HRG+Uic/uV0wUg9ryC2FyBF5ar/vTr
znZc1QPtXg3igtVFQpqR8uobByvIXWszmzDr+2y3713FYOI18P3WLHfu3kFGEiPm
f2Qy0abRldRCECPInZNZvLe+0MvJh2CyX2lWmaxrQQ2hxLWZWt5z2UGRU2AcojbR
41DeupZ9v3ex4OIQP31KixdhyewdaGeQCK9FnKWyE0Bm+Hi/pmiVAszILZQTCDN1
0EV6cPbr5EbRvFfVspzle6YSPUdh3prWUGsmYB7h8A/1iU7d7tbDI7yYQEFzQAVc
YH7fzxhmyNk6GhQUdnfIhjlusEJ/Zvfg3k86BphDmQphieKVhfRdkzXLUtVlHm6R
RqFiZO/dgEKyLo/i9q2OiW6e2BTrz25ULquERk0BJUbGEWCnT2O5KxmZW06IdNWx
iy0oxFVhaSKQxtufiHbpU99AsUOfzw8RGfKIJ3MeSOKXiMfcDUhdQFvBWr1Vi/lR
Tk4E4OGTHeUn1RJDQLc0lEN5htUBYp3qPAqleTDzh2MYwSdNMLhB4a3tUwANXf5Q
OGEDKu6emVxmwBJpWnWYJ/4kgoUywX0tQ6MVDBAEDAYBqEULV3NZBZBm4OGUFJts
kvgel1tJH0acXP8sdi4GEH/AqKhIrLT5qpvDhQLK94QgtImcdL6oUDI/zWJEmEoh
bB4jSGEbbxMG3dE9wRNSMfKMFnft11FIAi5ImuWL9Pp5P8pd+TT2EKq0GXXqTqm9
Zp4ZPbwyMBOqpngPMTOMfkRthqtSHyubsMwlMpKRaKaucWCQefyqJRE4OdFX75z3
rv2vPaTP/D8rNSSe1PnA6nkAI2ZXB9+PCRjAt5pVbIS29tKEBbppQVDCbLdbJ5vH
t+2wneluwwFZZtl6P1c09bm4Id7aPEAVwF+KU3HFS1wRXUzbg69PAeJCmYsFquci
UaSDNBPOmD9I2kZBe2bWkSNqBCLz7uFHj4F2/ImbtGI1+MpskUIv4n4jU+52ZYT+
itI2BO1h6LLslrFr18wlKIx/eZXi0TbQdfdc+BXfAzNVGtkBRcb/G5rOqxtXWrYW
qP2hS4KP/eUoIlkex9wL/PsRA3z930xbCxsZg/D0OsS42fAdnhdndKhHm+ZVKS/B
nQmqzFLdwOL3ibP7SfIof+hLE119pvP1vm1aRtKLBoIVQXlV6442dRe7xRco7NfE
MSYUZVMP6/6Yjydn/+JYtzGZNwh4onX7bF1/jD8YsZwX3L3DdgUv/u57BOE0PKrw
aPngEdNvfnsoqqX/ASJQaQHmFUA/GJ71WnascNEqn9yuyd8OOIVuaVTlH+v7D2hs
TV9TCFEi0irPdhcL5w9bFBbexJxkJB2RVImH1eQgQ7tbYtiGHHGVNC7nLBRcUlS1
dxLyfFmKDKtp1raZweSImA53XCgxK3l1WmK5YDf7BsGr/nLsHmv2wRDkF+cWO5qw
XaIkjkqAY7seOyROD4PxRdKTwFphmhznRKeznHDjzLcfh9rppYTOJ4XFAN7OlDes
Z/t8zd52hKi6ocxJbZfLC4T4ZhYrtny91+DKcCfyBSTwgRuC0giNLH8Qsx2fpyFo
mnRAGEJaXw8O05+SeFxxjfdnuM6AOlusSuxDlyj1dqfO4NxQPlfkSE3wTMWWlZL6
6kYrBsIjFdCYVhGsQdc8gmeKMtMy1f6bUt+AHt4H0UYdSL1qaZs/pUCFadmjpqAz
dd8IMiEXJv2miZNOHCswvTvZEudwjO3VqPThnOt4cclsF881TqbI83BXJHK98N9I
0T0ZHEL8pDgBkfOFPBOa3mPpRPb0JmS8dZA0wl3UTlxZJUvUyGLsUPu1HLq6DwtE
GxjA7tXC1mgqBtlTSU7RjytXhpvZ7K3cPF7Vbh7o0tlFO3gc/d+qtH66I/d7yywB
Kpn7rpis68BYkFNPX17pVZuEBIzCH9WenPHROS5V8jtLiHD48yK3mGjI0to47SLs
rxNS6WWsoUAM7bDEQl/i8TMDQPva17lW/LcqDHpmcnzcntdKeSqWMxqXIZ3iAahV
BCSAITyeBroXsPXvQVxd7Q31FOqow8K1biXe6+hBZ0T/g6dJcldrLJri0RjEWZ//
ZmLUEpXQbQ92FwZb0OkkTS/3hxQYzUbmJXFz/5IdX3khVf+X76nt8eXaGLBdh0on
8KoyuVNS1o+jBIipoHINooMl7B+NN6yehdHf2Z5dQAKeGb/7lyStSlemZS8nd7QZ
p/RljoR3vwq73jzTYHD7Necp1WReVfMkueVrEHrZAkEnkA3OZw2PzYp3NEYDnOKt
JcrGySj9oiPw0QmBkwso+/lhed7IyRejcFWhSDT/gmbZs0wJlWnyCo7KqoyYsjSA
9Y5s1JnhamZlTzlXsV2cSyc0osVhQPrE5scySeU0w6YohpegfEaMFVbwyJg66Y7J
w+j0AoGdV4Bp4OoDfglq4KpwjkPb1Y8/3ORj+rIy1jR/q/wKQNoZErKwNptQCz5b
awaziE8kSKhgasMopumWxgE/6KaKZBhWqxYjU+55dy92eVtH9k9f6GnF7YVJa43A
bOgq/nL6IN7nznVwu+G1YIugBNb14cLyFx0nzWpJ60Rjl+e/4MCCNgNDtPYdYWIk
PtSvFH9k4Iszx4IKKr858Z6HdGWQmlHGPdCjhlPbPjZOqhD4g15wPj5l/WpnQoUi
XsuG2KOVQOiMokD9H4n2lFhBDYbgP1HZBVoVh20Z8nVarLWkL4yqsu1/40x/7TAa
61jkdUgpBvw6hE9B5LvdW4KJNxXPwpdXSIkDlixy7MTDzMlh9/oqdmcZueIC+Dl6
c1yTG4xvn9f/M+9PdBv3miFMaecG+2OKv3Mr4s+Ukj4Ag2xnaOkpXBiTDre5IBAf
3hI3W2e5kYj/nXOVLwOU0J5KN9bL+/cRbfatfco1CgdEnIZq1TJIwY8Ib9YrjM7G
phRnIhKrVBOd9kJ+QyirYOsX+fcqL/+s1zzex7D+q3ny1EIRdzHbmU1Wuu8f6ViU
BUKrDkzBLYTUpirtxalWQD4S/oyFelUTuV26Bha/mTOPZYO3ZrMRTQzJbfbh1sU0
I44LaqVRwrUSmZNEkVu6W/K5m9Ue3Tc7v4+XnLgGJ9LLp1a0UTHXm/dkrd4lwM7U
5lLIIE5Q0nDkCC+CUYv0lnfxHEXZJKE4MUgtoLKgjnWlWG9uvFUAGmReIhaS6EMK
FgMcDozn6h26vu2yny+f8EcPfDQWBtdFE4sai+7M9L6y2Lx8fS7ggx3fMPvpBNSN
LtK/RsTqI3iEhzfFACzWXKQz2ZvwneyvKCoDX7oT02SPexbiGOEqLtBn/Ud6ku8S
epZN9bBuk2fuSnR2kw1jf/Y2etcc682vCkg4UvtQUzqbrZdI48yBYMRMrvC4hyqD
FeR8js9zWO4Tozns5oF/KBPO7X6h7THGwCPZXrtLCjlxExqm2NCRpcWnKIIBi3HF
Hdit4WTMpr/2Ba60nXPc6YkdB+qTyrR/8n/Vh/iB6hMKlOiJQ+wE8i5PLxRluR3F
7btGUqPC3xw2Z7YqEnimv44tD20TjfOTIRcV6oY07WQpKqCjJ3/yq4iqyfF43x6L
CUjCjvIOPjcnYUcGxfM32zorLP8pBRaGkI1o9JOZQsKsFSod5J/8WUVqAEHJDP1W
ljgmLB9BekdXoO4RYOqND7Blf+6YgNTSvl8sKen1ZhIbDfcea+2CE2+1i0o/8uVW
rNSWE9NCvjlyGL6KN5x7vAXOR6pK8KexQVOGmDqpWDjEyKgJY/Qf3Dso4Wj0JOWp
A8MCt9Ypxf3tF1TqfjGv4cN6IQI0+kBpKkfPxnDl5MGz9JlKQFWxs5H9Sf4Gcuj6
u6QoiKDJpHjPplEvuD80QNhEKN3KG/Vrwe0qnf5gkKAgJxjKwU4u0dHWglI52np1
jDOZOmakd7G7U/W55MYqyagYNC/KlfdfeNqzn6XI7QdItmQrhgFt13Hzwv7IB9nI
X+NJejZCAnCjHephmyqWnXXTFOaWxigKpN1BD5irnIbz9/rDcLVH0db/WcvDmFAz
RzNe/F6EoCibmRy5Z9PpXVZVZMqZocs6+zFfsgC2hY1/S8YhBPMQK3LelYrNXGn6
7fptvSo0Gsnb1GGVOc4KGt9bVGnYf0k5ZVjnFTIg097i49C2qSnkh9txwq8HJS5C
7Sk6F8nR2nfhMWhnkUeQZMh9D/gf66Dqpa+yPjuuVH31OaZsVxuhy3TLmQ18fVSB
EsizIGU5GKV5yFSl9nCwWtaDnGdMT1xJYS2NvcfaTQJjJGTxaQd6NhceutPVMCEM
abUulr4FMtAYJKfFImXBkzV2cDSyNMKOinBpUsWezzhyt6snBIcnjkiIED+zv7rd
m39kge4/VufWkjVtbpnuNkl6vbK8Jy+d5P4t2LivGmuENfHkeicqzLqf2lEAxsJD
liQ8r208w9d5i39qF/UGwtloICvNzASLxNpwLMtru9lUcoCOJ3IFhY6wCSMYfuWP
nrU3/MxJm7vJR5J6wevirmL3i7LpXZ6mMrlKiDB5l68InWn4vurbv0iCCsy85N/y
ac5M0is/RoEODMoOCzFFYN48WelcOoylm1SA9Fwzj2HwkEVxjFR3GKbVAaA6w4k9
/XttT8pYdHE0PRZShEA9KzirmnuX0qB/a71cDvOZE5FzK/Vh2hs7U6sQ+Igy94mJ
F4zB0if7KDW3T/ClpuRuy7eltX3zCGBIRqVEMhmtB/xZ5hRqpmfVPxHDbn5KjUW/
IWwpBQbX0rmC6zPG3Z6oezo0YseAw5BSFTBsyFojEPREOAZG4aAW5wA0c6wqiluw
0QnkwfGaKeBnI3kRjDb9J400+hxhf6zwjXTkyNDPhcrkclfO+0jSRR3ysiOlboNr
m/6Jurb9w0C2PY7oixifvbpYPLTFFUXd/02cLm10zTZ8kDnFoE+vbb9PZYK7lDKT
y0FNZTTL62mPzBwLV2nzRBaZtTyUtkUNPPKq+5JOr4jS+nM2Gg7JbKnE2XkXHIhG
b/83JTV6ejuLsUfKrNXxS3NF2jnSv27gLeXMTWz02jPzsQtfE95T31g439AnCeUt
CTdhVPaGW7ZAbtqngNbo0VjAzRO4TU5Cnn4F5wRYUAEQGB6TgNv5MEVMrIM85WTr
YjaKXnyyPhLWN51zCiHKZVUPAws76Gm0BpPWFi++nd/0Kz/lfEMCrNTjl14ZlErg
jSFS76nqDE9H5+dX4CkOsp9GI4joZgMxO5xat7zmy42DCOXi70LAVEfi0y4XxhOl
yAoshP9t/NFWihj6MDr2b7YiBA4qdJ2Ye/jfE/tbf3KRbxDoe+/NRkGX8MX51pQK
Jo7B24hSjnN2gRpgFbrhhi38hqby1CAFPSAVWl2BXh3dL8EgC/HjoWtm1vkzeFBl
deykJm4KDu2Rnby5uL+Q63liQz87EXA1eImkEzkvKnFtpKH1+RHZXl2DrkQPWRpa
qI+gtIiN9d4PGLyXCJUnunfECSWgB6PYudRIRtqf8WiMLeu9SxWjO2mA55rtE5L+
MtMjgOwiEVvrMkgnJnQAkrKfNQoEmFbi/l3L2cxAoW94oSuuMXPbdNDvjiWFOEei
5EVHF7Ij74ivu0VHhNBzzvVX3eBwXg/RhYA26avqHO1GpY1Qqy1vBJOcbFbgGitZ
HdSDCT1cTzNPVgviYNlqQvFcT/FcwQuy4Mfv7YOZtA1cTBAdpY5WdC5x45VDBe2V
ppJ+8cXc0nHaOAAhIkqBubb3/uYagOGwue+kSKz2+QfjD6R2xmQfkI2tJMsSfr1K
Quo80NOFNAI2hhyi2AwYoAYADTvo6yLrJ4ZvTDlRelcZUIkvr0+vdGvNP6xmfHkp
HQtV+KDXZPQ1Qw5QEy0zjZ5lVH23ZO8aocVVEOKqshWfaDt9doeNYMy5jkXWZWPk
TUlDJEvgmo4Pt2Bh5QkKBzrnaLDTvFI97/FYp+qbxKuhpppcOyDZB/mnBk1MbbTG
Imo5S72+r2BCvSbojeJ0Wq0hc6TMP1ZaxlQZxoIbw7AtmzxZSdlRQMfNGYpkA3/0
dACAQxL4gBqCfduK/GOKURnNWOlulMFTzzk/BobKenPzyp88kEZ1SMvfvxFzU5th
2i5KC9nU9zKDKAWIR0dBAAlPWlY68PbQlsyqvp+EDGezI3YIo3QoSdjMA4e4FuXS
SPIibc0+sijTvLvkxbEwu2m0BzvjCthJAx6J3btE9OQ6sFrZm3ZHKLWuNFWA1QPB
CcvHo3R/F9g7AqmCIqNI42dPHCpnZLfp1NwBzyVfgFrnR2I+YUU4dMVmUC/cON43
guN+PLRPIcpEzqttKhTEQG/ZoFeqRPYUkAJoWnntL1vWeyCMdEff0x8leuQu95od
mZKT2kOxbhGTnwcvyHDnGdhw1uXf8TIoyuUiW56+VgCpe8b4ujetnATyVy9viz1Z
eO9v7DAFu2Jn0c7DW1UdAdl9I9uGPNFjSEhf5mKVHurnEi1pHzPbzEvOl7R/Zoje
LgCuZzlrNb5kbnVfMfanlMWY78h9JlDLPutHilEUqnh0HTcYBz2q7K6+NW0sOyL9
4E3kAybnAXDdZf/L0q/lVUw5249/z8judGftfgYYX5Ayh5MnStjGREdMGBYWk38i
YBUdq/1uTbOuI1mjfXeCPvvjxWAL2k4eh7S6i2RaTzZDSOXU2Paj6EzkxGWD76B6
UcMbkJwOCfySf/cKZlooDqSPt58F8GTboomxzq8r2FqYkBirlcD5VbxZOLUA+OdF
R/sIJJtmrLH0dxosU11PwzqKx5h3PCkGxv64UhpLMNol3EOapS1zsskP/6KpAjbw
t3StnhwP6DZzC5Ac4lsGpO3kgdkjX5jtEecOovm2KIPEN68fIzBLyc6yf3DmpEtf
H8nSsXkif7kqQ1RCCzuF1+mQadql9Cy/T49tn8E3FzOIbJczQQJVb+h2LHwBwezK
LyMP2Mue+6qVgVtpBKhZHD6ElS5MrnDn9+JTOcvzTJ82WrTqIxCP50LJTYO5ppPv
5Fmm/1z4bmjan8wWWnP0IQbW/QsYK/bVp6GBFdwcHIeIGRApZAv+o++sGtGkN9gp
Ix408df/Fi+Mxpb8Q4ECI7RULaBEBfCS7+uC6NsEJLqFpqyp7WsXug7SOZYLtpWQ
+tW+LRpiBgb9rfKov02gYiO0ArCr6XOHlzPsBo5m30SsC7AuAVSFcfAPoL4gBKOt
QE4pwQfW+i1j3283tPp9TLBG0FdgWhg2o2SD8AE3jLUzAQBQcW5AKFgd4Y8dozwg
7atEGwe126N26Z/q3SnmdvYCKEATwb4Ks0ZaK6fb6QxwiefH59TR78eHb3ekKhly
L02dYT+fS2KmlqMACaHJcghX5tW98AgkBR0zpXGgbi2WjvNLM1arrDdSil7Nwu7Q
ZGNhuVaFPf/q4XxoR0H0B1kwk67wreCjm30KfJdyebcuiUN6t1EY1D7PzQKBIWML
BmwGSey6SIX69IzGq1xHk2e3RVXQtSva+qi9B+eBuVqaFgVSA6JAvxyjhMANI8O6
TQ5sJ75gTk2FztNqAReCbgCExXlwncJOmC6JT3zlhHzcfl63Nxgd7xa8RZq145+Y
Bx7XIWKHgU0D2NC5zREj9WcuhYk9XD6/x12F33aDnMxuONBh59MovMIevBojByCp
syaJnz0Xi9C1dxMXLG8OeuKFUak9vmiNeLbtsEEj6RqNcTcaPkmrWf1cjn8zqX63
+kZUbMyruoPcNgf1ZaYZAUgPhGGjpcLwz1LTcDdxp+xQdYb67OP1R+cNEtgMymKI
ONVVsYATxdD8cflfSczLP6rX8WzcwTEgucpIOHODGoTVMxRR5+yfwcdSZ0fQIJFt
aN1ItzKk42OAgfzYAOPwApoTJ4PSHVYojRmlDyQxdUA7TYu4Dj6M2/ajdJpAIm0w
gFGNtpof8/zvFmdfRXSlLxV/LSxkPNa70El9D9zw/XTPsLJRJWYJS6wLqk2G6E8g
s5XnlbOYGo8ijy+3sRXyDL6YS/NXdDLmrX13Zia8EZTgngWtFBvSxNiAK0D8OM5W
ukIbhub+JQiBQsC3ajGx6H3Ii7URACcwrdtRVPe6anhNDtscEvQnODxt3fx5XQ6B
qEF3vsHxoMospfij64gRw0PTVngZUan5poNnVmqp37qYklObWVqylykFPPIBfMW5
x/IF7sdaUCzF58h37rfto8Bk0TZyWpjiED8CzfIg4YrD5qzlgzBCD8k4OMN/5H3q
z8IXUquhy5cLlneaW/vvF1fIrmPw6XuayyELvgRY/uW6+c++q2t5xqzbUHCBPFSF
KZ//fhAG3Xl9Lvw1tLW3hbUSpqKuRJTXGucuW+C5ENENDInjYQLFufjOhN+LeW8b
tW/xjK4VlPC7Kd5tiBLSJr5euxqwJiVmY11Mp4widdmArQiaUqueMMGDawIGgr/m
byVuTpPVhycWDvcZRViN/NU6DXtlUUecGoDS+8+eJr8vX33WeouU7euoCQr11mQi
YF7/MeDVL5bNpKyGn51p8pqax+yRo733EGu/UaBpnRDP/1myFH6pveXRyuF96SjC
P4YGYnTO2I0Q/huRuNbfENoACJGmvirMuliX1kXjLBD5gqtOiDvlOzlDC5x0F28P
lS+kNVdudu2x5XztTE0r940pgojpTOxZXa+efAPh3Y9jLUkS1y6fkCRsWDN5xx2E
t2E6aHCSA0y5S1ta4/nSlWMattI1EP61M8IcBuN/Lt3/CNK+kIh6fwf8GaA8F2Mz
vbFTJcbulk3PG4L7S/NJvpgg80bI7Owvs2fNIcIYnWwH7fGCDk1dpF5tevS8FT5k
QsNBaxgvhqMGAieUSidJiZQkN9lgu+qSGiJwZT+O3Fzv/vk0IgXOA0yTe6E1+NVs
iv1kQuVzU/0BJ33AR/D3biBxOXUOQTHaZDwFdi3lm0KwM5oqG9frLI8ysFeERygA
DTatWgOT4DjZgVDCTfjPo2+myyb9uQ81Tk1JZZQs9z+5s/Pi1yc4pcFCejF8tYJp
/mJ0dRNDEw8dxWu4C+kVDlVnbwG5y3d0ktasR9StjKzDMbzptp2q2J0CA8Oypyu+
zoklkXz37N3bhWslrp4yM+MPSA86R/4cDPSmtDDmgJQ6bG6tkMw5T9AzRh4JTmZy
O6AY07To/iPKHZVddWur8u5uraK6XpR+tE6I+eobFdq6ow17KsTedSiyu1EKgwpM
SigOL1jMdftA/vgRLAvviKMbs9XdpCvyHtLNbXajogZAItqz8qeVdCcPniAnIgCJ
c5FESEdZniFCSWtIsDSNg/hydliSJJZAmKnh1oO0ESn4bXYZdKSUWq2QlVBMZwHv
UbnMbXcSFraA9RBIMy7a+VtCaRLx6FHxHjdW1cXIeWsYjIELL+tDahsRiOCm9V9f
KXiccnHScpFY9PX/FarGzy18atV6IR38AQa1LjtKZhGUPk0OQlzqSC4+546bWS+W
+YlWfNP6KHgxwLbqsZuYebuP1VkCVL0bo3zeW6Ydqd9H+7AGeoZ5h6DrDpfYeFEp
X8LyQvvDXXEBIJ76h/hUm28usSOP8Ae1FUwLXJsd4CrVBxkM4/0XNyBmV1dEFLeE
Pk9qiP5rwKo843fnmMy9DhRxvLFkhzqGW+s4X4LbWQqkKftWcdeLfaeGO9oGU+RH
0XO3f3pLBijxZS9IvZxfKEmVKg6N3EjjRs0PtwlS8rxwOKbq7lFVp+Ote6hiEUls
9t2bQrNIY6f2WzKGz83KDXdgHXwT2V9LXdiZJAzpESoPsJFvjgtUynENEpAtCQlk
jNqy7a2D6dpRg7B98SNiyOf016bwpWUdFHqSXgWhLVfdf0FnaE79o+dl9DQpWQz8
XwD7ORzjJxeDKZ0K7sZDG6a38JOIOi/b8Oo4CKQgwZkZMViU2X7SrLmLZvlRUP2K
uinWPjLeCQCkJ4dKELapGiPrHK7NxKfcOHrkhDgQgDqkLJfbjDgdWBbb69iQklFb
H93lwAue8soiW+OF8vkwHiTi9BziqS9AB6mc9U0YEkOaqjiPw7SaOSowfbqpaLop
4uHcsO06Ap1KyrvhmI6zPCGAqDxyAD5Vmqf+D16vNQVX7e5QSfQXXvOe0j3+b14v
IFLjRLc/33oFqsjDRHV74RH+VAzCE6wUCkuG/+S/euY8+VXbyXZsAANj6E6LXCJc
QH3zlbwaCzjDz4hSJbCH9w/kuqvNe1SGwxPf2Y7irZG0GPS3+d/FMpbeAezGN9nx
U3VHVXENIuQh9xo7pTKWUKBbc4lv862THFTx+Qi/l3BrJq5GsUirbeWaT1N94bAh
rARxaiBEskvOzCNLfN5K/t53VIjvPD8Yhhw3XqGe45RWwGmGi8G3p5bhtYPy63wb
08RbjQf/FZ9hAoe5eLCacPpMIIEQIviMjlhy6nlGy/U4uPXCxv364lQ5pJE+x2JX
dPRIwV6U4Kmo3j6Fd1f/7OgTBk7NIHK1OENlo/bGrwNObzzuUvtJiEepwn8qINOf
a54VvM+IuTX5IMPSx4HaHs5T+/WNzQdCNtxXmm/0CcdJRGR5bm98+Jidaq1kIxcR
QMt7n31fpQbOwf6qvcc5JC7rM+OhhPoCgX6zhVugBlnTkD1CCerUXHwSd+NPZbBv
p0S4hB1BcPIdXO4r1GJX/gs6I6diHXns54LsLA66px4xIcYD5L9ynEXuIgSPHxTz
juO1Kj0K6BbRC6KVqUaxxAkl8udiIwcau/I+hqLWy6pC75Klb615yK5HVCLngG1I
ex7XCJ3gDGEETQR7+0aYrvu9EEiU6tWEN1GPiApLt0WJpDpvftQLKdIXhnvfVe1k
lUnj9yz6/EaXijxZ0FsC7Sk3DyBwek2LHhTxyuy5JqJzJqt7CsHOkGSLc5X6khtn
2IiGZH487PyWnteORjUxLdNzko2pEEYoyzV3IElHT6txaLtjJA5lvRPZBT/J4Uuj
8CcOge9qxRiSFWF3JlIXuj9juxYTUVaxVCeljuUFJebTdRC9zQO0C0rRm7oicqt1
FgPYAR6rop11y8rGDryoAS87Gzh7D47yki4RBwFY83DnPHMYCK0kjvo9U/TdAQzY
gVKLrMII3vIpAmT5iZKUq6rbjdSUBuC+Y+9XoLYr6eXdX6EdL9RtD68hE4ML1vrz
A1Hn4z2O5P+wf2dT71XWvAIj7eSCZ0tKPX1Pov1gaf6b8CZpsPHjR2tRJGj6AIal
NqsaUPO3thtG2d9NKIpAjcmkuVlkXuCtn9PEa8bmcVvUPvP4sR0i64idtDOxJQpH
cNqYOFLB59yVmvaxs4c25bFurY7cxO7gGImqR2ZzOzRCz5eFvQunXDDaZBaxxicC
1ZDipoQFrWu40ChUdbUJ7ihr6EvEn6W7RDAQiMFCsiZ+zM1pe2V9mFooMTBWbr5D
exbAy/9i3XoeJRrOaC+ZUMMmerPIimKWJngos9si9htuY6WE4KrxQCrlB177Kt2x
FPjJ9hrOI6fb/VstJOskem8H3WBT9PZciTkFISwwK3Qa++9OvbHWc9bKeFh1+fx2
Karknnz1/C29CkfySyAiqPdxpIhSpqyy1eJfQPROUL+EvUvinxV/BtdiqUBHrFWd
YgM8iVDD08lv6wZCt4u2qKfgdECXQS/5VpqM0DGIl1Swvtw1b8pmhfbVPoECEoGY
hvFITXCiSaz5tL6CqCU9yzmB80VwiypqObigp9FIQ4lVseJm+fm8VptHer7vxCKU
U+j7zoQ0iPs1lNXa8Pv5ggjR2661QT2R9UUB5WkVgA9MMFvcZrMS797/Zrd3YNsL
nRQ8iPouusati9g0+iZFIer/b6TJL+GjnmNbV1pcpNNgrdmx+VwJFJdSNYwJcwUf
TioXZZ3So/FPiPRkqk+p1aJRcLzPEsomz0UzdZc+eT86tC4tvetENequbnqlojqn
BBY4PuwBrjnsmZpBfIflnVLtXKoJ5PayWs31MxoLJr0CnPosZ+jwrHbUXFipzW77
0ZmLLD71gdaqbJg7PM+xN6kPGBSrK2ss6DKglSvK+5TSaLsD35Kyb/V4+HqyzBwk
eNWZ1L5ltV4W8adC4i+PCEGmjaBFD+wvOewfzmJwb7D4C91kb6X8tNr6BzgyZUJD
ypJzU7GnJNa/DXaUe/VXroq44fmQjEmObihvMtfJIRfR87Pox6H1+SP/3EDRE+WA
LdBTysINPgENTcXyl7JBEVniP0p3HuJtqtYmr/gFesfgrJrjBVTTY2OL+w57aYbY
K137Y+ryZzndVYNOv9kZTcHWfFBWme4O7GegmSI39TLY30d9Y/trZegdZWWbY6/g
5ok6M72Vpykl3urZ8F4LIAMWRSKLlL1LgBjcSTko1CvJIB0AhEo5rV0K5VRZ7AoT
ipsiPPTD94ZDX2+vVM3qdeadKYreX/NM42wbiWkC+DOXk2nXB3Rcsqbu/AjNudym
lQ+Uip4xZu8L5tzIJaJdh8tC+yTSIkvBbNQwmkTpF/lyRjWDpKmboGowkdMhvl5T
jN5Nmb1aAIhcZ25tN3FnAu8yaVYuY/UbtClMZNtt+wcJ+x7k6sfBmF3OKGkafMCI
LAjGJzrA7booeAMgzt3zHG2ZPK3wdgBKSGYdB3fqhL2wpgTGDo/CpuPtDov1I/x5
/rNn/6LN/mdytpIji7FxfdlpHpiN44UuE2rXaj1tEuGFz7uu+kjvL9scGVjwl7Ls
l77fm61MpoGWjCBEiYfl+hu58yddEwUwE7F9sBFFC4tGuBInWnka+Y9lYELL6AeQ
Ff4RBBGzvJU08zHTk80EiZRpOmyDQE5ZEq77pwVmLrxhTKE6mFIyc1DaacZ2QYsq
OnLiR4Hv6n2ENAh+y0X04PGlEcH2FDl5Exa0Q/KTXQ7nR/sEhVR9SULExuUP7fM4
g3Uu4HnyzV/TyuUJs5yOAAX68lam7Y+wdk2UxIb+k8Xi1eqIUtscWyC68/OsdgXI
5eRcVZ34KJkmKND+SmCpIPOB5+BaKRp3GfsAgq6DWYEdk2SgkTVNAPvVSncgXrOO
C5DyoxCtubO+D7dUkSnRK0d7YkyLWBWpmKPqWco5IQ27WKtgf1MCe4kuOfcDTQNx
vNOrMozd9aDBdvfSFJIcTLsMvYN+CqlsjSiAUsL+y7D0ttxWMCAepc6eU0yjrN/A
UCnP8kk3gPv38y/KNQsSymTTa/nxCbeBFyxSAmhJad18Ai5wefAnnePnYHyHHw2z
IT3AQHRJHR8CTK4OonXCrQzVD4pefKESZk1Ypa6pHMRI6dwKU7HFaxJ4rTFmcXjP
BTIv5hvEj08SZOLRdl+bncY+bECy4i6dtS8VdAoV3VkPJhp0p69eBIRE9c9G+8B6
HlpSZM67d7yGf4J89pmJL48r4cuixBi2xgTkJnj4CoLkq0g+PqDYIRHN3uc+Wrip
sG08SnsbPbKsucJYzSa1wJtCGQS5LQWHa3MVbPGbCFTTbq6hWF+cSIMGEcHmrfxJ
LdgCL6IQsM6XC8Hl6qwluF+H+EnvHrzu9r4bxJK5zajYJMTkJFWtcuhoGdZZi14r
gpRQGNhyYZn49L2U/Z02ViEzZ4Jj/LZr8R60e4XjXolXy1eBJV3xzJGNzoR9KyG3
KGO/hD140j1c8cng0399K1rva+i9RiPDj+k0yxajDBtlZNsY0ueiQDb2tjb+p4ds
LuUISMseVybGJJb33akyGvW/q/TnE+zvXai77uzzdAEs5Hf56x12I80OFMyWcioZ
/B26bvMa4RXSvn+yegGWN3TsnWv2+0W/A/G/SzXhMOzUk2IF/2LXq/cA2rSINvlo
62WJyNf1NXqdjhXYeYoJTXAPZFG1WSmLWTNGHX6d/1krdtCioTNBCGYO1annp+Vx
bDEttmN4hgWffjieg/OWjnuEruSS3huspGRg7hHlCw6pZi8MOnQPpDz8G6ECrPG6
BgWJ0bt5fzDm0+EwSmDz9L6794oGdVv3cxyCObwNAxsNTmN0j7j0l4EDK3BmOSEH
QbHHXBLugTLEGA+l4g/Fzm+WE+cdYluUEnfugdZWrCS1VUU+J1/EnUBXNL+v78OC
CEUTmtCa3v6g98X7gFTlWF8hxyJzI9hDmdHLCrZQzanwgy0ut2Y0FuLthfZpmzE2
Bugwf/x2ROjCBEddgDU10LOiVV0oFoIiA3/7cGe1VooRwsk+qQJWmoUCf7DyFpCb
T/ZoLaEANr0N9OKesTxEd/h/ePV/2w3yB4oSSj3xvbY31HWWMyHoGKKtVp1YY9GP
Eg8ajEZyeBdmF0Jqky5GC7wU3rrs7Gf0YCuvOqg01xyyTJQSXMHTRlwWsmKELKk6
iN42RBJ5dECXrpJJZDG8xkREo76UNExxsgI5y/1/wGsHqmgobw0X2OSMA8lQPGMD
vTTAV6IPIbC77GzGZ6toobsvGTCqnTYfXHU7kqyECfqnK/97WMyiYWvpKRX8pegF
tvauSQcCPyehUZ4oTw5IiI4XE3UfjkC5CZkDrCRKkM7Cex8zBAMIeHpUBsP6i8js
mjPQI8L6Lm8EhPP3QIdb/46GPMkS4fjGX/0yWCjZi1s+I8lo5hjldEBis3LFv/FW
SBr9DDLnRLBM4WVUCsMsUZ7WRFKIblQAkkLNT8sPHj5f03YghQGaV0Pcyl8wTJ7u
QXMkLqdmpCCBVtWnLqXZb4PetV+KPEMugP/H9vr70ASRzpbxwiojHZVuX0VsAMZp
tiWn53Izzla0bzWN4r8wW3NH6RWMNZ9OTAdILqkgC3K786GE6Ihj5WvuN0Brhlyg
shILD0gFznDoI6v7MwA2zI8b4N6K4mbxK2g9/zKhmUlgtJJPyUzCNwsQLphoGZq2
ArEmbBOsmO02AdXP/exygnMW8MzYvUSGgqzg+IkFIIy+0HL/P+d9IQTjm35iHT2D
H5+g5TO648rAlIc+RxvcrT91TsCn7H1esNzSiHYswbfxCEXxfrHcgO25xUAnUXAt
+ZPGnAgU85AlNvHLf0XN/TbgKX1cfBCkRxHcim7LvTbe+KnPTCKpbyDngqXVbffv
OxghlgLwJ5B+dee/KqOTivVfooYgxJHaKWKIfXERGMBqyG7vS78AYKyBF5y7xQGQ
H0HSOtsxwEa7OO+hZDRzDXU27rW4o0WyBepgpaDkEaJl9+WOZbHumAo10eyP+kff
IIiwQLig4f0DOJHk/MFM1rNoQYJ34/ELPFAsJDXr/bjD3UeHLzEByW81sPBGCHR6
4cXIph5B/8EnCWoMJzircq30KsNIfolKDvd4WU9O5DQozAQo6rMh6yrCoPZ2xpek
QRURScZftrqoQCBVTq12ZWJvJtWaeCgpjDP9tuykAhfbqHyF3rvynnpQ6VefL7G8
7K4w8QauA27y9MeIq20Ua9FduDfisfJJxioNtw2J3KAsKrJpZJ2dtwdDw6qVFmPs
kAPshZkbEhAeb8KcA3gEVmwmze7t2/V8g/5DGg/IedFmy8hjhik3p3hB7lfcHBkf
zlMjKEKb+X7qDoLCfP3NQ18BiynEQIPCeK6pI8e76a5vszUurLXgoTkyYiKCEmoi
MoOWFslfy2G1WrG2ST6hBPZtlplvWbXdzmSvR0KPaEkiBBrsKaOpsG6FDs9ZUQSM
r26wV6PR9CMrInc0NoLZzvZRB4Mxeh1QrypiDIVfBTVZJRIPu8LLm2JN8v42paWW
gBZzBCyj9uCUme3/8aj2rlqXQfCxZ8blbqsf6/RQIuZxdBRNeL57/91Kj/o3CcJL
oND2j7+cMoF5zAndgZK1/N1t+jKdpxBWw+AZIu+ZBobfrNorRAa+4QgZ5vxk32KU
OOZ8GxaUBEatBKnYKzVbAQHDntucUNShZKtzHBFtHcMVhjN0weKQBcIhybIipCkM
QCb7FpcpjR/HAL50KOYvr1K6sj0UDQkjBWnoYvNJdrgD6p+U8aZbYTqJBowx+liD
K2TovUJ/qdRc1qMrkveVGFGu/TYQVBo/zGTJfONjaRWZulXmS1cJ0ZEbyFr3vWSJ
85c+xgeCsvAwrymF2QanvZwrNztLUmzVx4Pn60bvZG7lAPkQV0ZfsPuRj4Dghdu6
ACRy01Moy3JA3oSrPW+3DMZavvTuexcsQ7nECI6u1yoxCMTB/y7r9AsQyBsC8GaY
f2tvubkfEdlfAL0xfzoAJm7si1aONEK5bqZrP3alBKQDYEBXu+vd9mhHktoWW+Ft
YT3j74IJjmieNwLoFG3+m/9CkbHXriGKcz5uryasL07OGVcpTZB/ZvtlIaHn8rag
gzaUaI+Nd4dSTIRLUHIYN3tbEXESI2uXhaNKOOirTyOybKImcKhT1j9EU0h/e6ZE
wJfkKmwHvHV8qhYVKfr0ppdG3NhMdAh1wLYIKTDnalXQ8iPiKDAAjvjRv7kcgVFi
2343+KoTxe6qU7+fjeD4RQtQrHYsjG5pYidwFY4iCTix9qaTLiuvAKJVL+ZnOohX
wbsHs94Tw88i8cWPrH0ZDjohC7h5z4q29cOEdwXsIGoqmUBFmJkC3/q/ZlHoQHTb
1Y9Oz2cvqWgVZlPqqHMgv6Kz2MysIKLPXe/Rf9Eto+/+YtvzRIAy8EBTz5hHv2ND
z30ohgwYBUoOdhvqvFa8BQVE+cYa/ytlh9VhdSY2ZEPy6O8gJU8k/9NRQSCx4L/y
2Wbd9xTGy+w1/f0Xf8xWLg86MQL58ME1KnTRca+yl4L7eMvU72FQUB4UEVxnd2TW
Tse6bXNXLFDRQv4/NesGql417aOmAqgFsPWBed9IH9qGotYyffNowvKQTXk/BUS2
zcNZVp0/lyqXcEDTZPDw5oFk7YuwP/ePdqrhkQwQrLPBPYbI0wrurno5EAIZuOKg
J0LWdsCreQgmdHBbIpGlO6hXUivqXEj0h3E4phgWDp27Jq8tgIcfJzW7KsVsYDvm
aeVGCLUfYgtxnRmXTVAANBzsaj0I+JXWkfZ8ArxMs8zBp4y3Aqy3+Bf6yMMtiJyR
YKoAyQat624Q/UMQgxx2WeHFX6Rr+odFTBpNmBpttsp9zPUI+zGMtuDB5HcZx7z4
E/6iMN9qEPxNh4VhAJtqqJWciTLugIEa1uLCjr0TjDDJ5B5zrK0pajHUl/ZVAfR2
RVAip547I6G/yqpJ/uGApClHSZNjtHUiwXJDQQ+VKbnVy6Zw1jC1MAcdEFxm9W41
0jfkdIdnK+D/NMSaJJ0NJEu7wsCnqP8e6/fK+YXwQe7G3rEFaUzAsVatnaq01l9Q
2fwYO1XgXvKSqMERxqxaJ62xQCmE6MMOnfGZQhLtnbBXbqmF8NaPoxqkJdiuLAHJ
WCeQxDkwjtvbaBgqJHlrEjg7cukJElVuaPhfLLQHClHPHeFgKnjT0xDZg1Atu6KR
OQIN5emAqC/pz1czpvdDftfnzmMZnnl4iDyuHukEeK7d4dxse4JBAMdq5QyuGPib
8O9mTAZ2bKD1JY8znkSpBy+/97oRcuFOnCeBc8DfGTO3IHn7XuGYUKde0RasTeUk
2EXao7im+nou7qLUAe+EYFkMnqd4wFZ+AoIsmkUQ0LARetGW2DMwtzDrNScJhMhB
e/Edx6ThkPtx77jeZplcpqmgH9ghpqlz3YmzlcO5JdSP9Oym06BS+lXy0A5ew0IC
e4lh3aZ4YAjII2NQAJiJAyCXAM7RYKKineLZb4hBejZz5xZgxpNj7MreOk0UkUrq
8LjgCKNJSKlDp9jr1aXyFHBN+KS9sEvHRrcCIx0+OH6Ch/VECLHB2LUGrY7WTWfj
DuL6s4XQUq3ZNu8zil2wAeBDebkkWiZEPBdMlAvHSj7hE4IkOdKtiVwC4oAdu0FP
S7qyPrp8AXpnXnRgCSR4Ohg0fun8mALLAEUGyM/kfgeFAgNMLMCfEbQLMPUhB+i6
PHKXrbAwu8Ax9y+W+BP2RXjBXm9lqZhLs5rhg0aon9/18AcPnUBtzWcAS45CpWBA
m/VrcNVAliNM+CWwiyypRNOXKM/NN4smeBbqXS1LeRvh6yku4cMAnEdnPVrlJL/E
rGqrlha3IArPL26KFd70zNbMrWyk57y7QaIZ5/c4QGarpR2ANGAf78nDZ/i1m+ji
ejR7YnLZQ43ZX3fxhLFuQQzNCEpek8fjWPaOugLGPhifxHdH1w0IeHjTz7ZrZyMJ
6SzPpfHSvTst9rBhI+V0wUQxLaB2GqfdfGD0BSp3YjaD6S6ypB1yHrBdbqHIltw7
zh6CCtuLUGoXO2cCR4BAoJGkjYO6cLaCgXQrRQyiQIjRR2yyHXhllO6h36u0UqEI
eF/EsQZ+YMZnYk3l/VdMp/XX4ga13d2oeoCajJKcdyJ/7q0DmkInBN9DYQe5rFnk
HejZDgphMlIE2l1+js/Ci3NxT86Ua1awAlbevloIg4aAprBGbTbmYj2dAVoOJrAj
1IJCN1vaxeZSSg+slLYwXTCUnV3WIK6xFNbMyptS7yDZ34k0jWGWGahK38ivWZOT
GGCDpFAv+yROzyJkpyN+bBpT/Lm1Pr4HB3l+bgrek16CdYQWSNN2CZacf16L/tFI
Cb4un74S3LHva4c1UNRGkDNOSoG2apLM4BqoKpzsnbFYgjLTPC/UTZwEFK7KtaUU
D/zSNhhCRp/YgG+T///v7+mltVJIkdkCl1JEpsV94fBP2j5H76i9VZ4SI0SY/zRB
C5BVkS8uJDONlqLmnXLYuTobxI00j3u3hcum+BAWJOwMSP56qfsR80Fzmbcenq6o
bcZO1c8Er9RD/jh1S2PvsilEb2gx7WXTHL/MFb5qbPQHU7W9CWQDiNdYAVrS8nAq
uZAkaQYt2mAu0K9U0BuVTteSEf/j4VyuCkLN5tnwrfUBQiR2ocJ/2SJsImWrbdN1
VwgrzAw9EZ+IifiTzjlwCOzykrExAPimbIS1WhYxAK66QuYghj2Ls4Yj6h4PGPF1
FLcw4WPoOdiqOkGv+ruw7P1Lfu5j+ye6w/l5MfUT/W800n2yBc6aPo+iFHH5WYmO
NKPaPlSQSfNCz62jJ/3SuZRTXfDNvpMUQI21ZPQpoe/zcKy1ZCWArdYH+Faa0JjS
8u2MUvzIp1xJyXhGgbVxt38QzwaxoXk/7o7Ub55t7uDFsSkaRDET9xxPLqgxsg5p
ah9HGXAt2GEiEpjQC4ExWIPOwMWQfW12ma78XC3zVdjt/3FDoLKbJx5iYhZhW5nl
1+oUeowo3xsBVAQhk4gkFyrt9i3OeiTsU0xBqloWbfeM7srSjlciQ80fwPdaGL9M
6N4adeYP3KzmTVjStzEbPE1fKUxpXjsGd6lUvVZAjGrhc3O4bFQoVJhyBVLrmrSC
9Ih2nWr3czY9UtCvYltRA6A7/GBvbjMr/VLalLhaE+3IFP/wN1fUwaBsKFa8aDME
qrurXTQx8Hz0YBWhfCbuq2jHT2oTVpz69glzy087bafZNBEHjDEY0aXdnJHQeFIT
aj2lFKLwXFLYFqC681c7gG2iQ1l71dx43Ez63qKXowgWMevvu9oVZFh8UfR2vX9F
DWcdU9cy1Ch5u1hKrnsBaU3J5eh+UAWYdl93JGfuCN2WF58CHGIfpzKgnA3KHCb6
V7C/MZUwGopHnSIpcqa3uWDZzuUReCQGza5NlX2JMt619Rs2A2fFZRNi4ZteQEkg
qE3aOmRzqjVeVt64RqsQ9wjBqk1sv+qqgdcr9DXc6G9yvOZS+5SCeDOg3/Kl1hjA
9TSL/Ot3lZnxwSAamBPW6x+hjh0SHlHOM6aoBUjrvs12kQ+UTzSPl23uF5jpOTO6
iJHEr4RFjG5iW/34Zt+QzA8ooHLlSVBHKxEh4fJtLPsbAAcb+H9xMwKLibouDXPb
RncWJeWXDPk1Z4tEvSssmckkuy/es+Nk9zLMdvhnYN0u/bo9KxbYrBPQgjZddg4d
hxTBW8p1PFp/w4E/xqsoNkxnOIoPa5otTQjfGqJHWXaZmp/0A3UiarbqSyT9MYde
BU+jrNMeD9P7YXfNqtqGak9HYC07EhZdpq8wrXLsw+2cSku35qdUvv409w8SBy6w
ToHrf5aFawD3KlKarnfpz+uvrGQFdAHzeaU9t6xwf47PKzBYrq1+EVGpR4t12c3U
FgBj5FBlkP6DGuOrt34csRpApf3FNH48ISBMeDrEzOj31CAXHo4PEPicIG7ieNr4
lEFzABlkShIjWJKzaaWotr3QaFm2NwAX8rW/GBghsfmRg7dhct3eOLVYyXYCIR1R
xibaYlM90K7NZ9+BL2K7FY1fp+58iA7lMmZGvW9u7RQ2LWyxO42FNU/6wEbvwlm4
nG9Vxhpr+UL+q0/oqp3/SRMJQaR0Y5Jj5eIfCYCR31iKzsOQpiV49bO+IGkcc9+z
ucGBVwGjj0wfp9U77OoplNJdGiJQBt/sVB8zI2ycGocszIP9TW9uVgpD1KGTevH6
DTQrNWcuWcLXLzzh2wL7VyxJpfiOu9e3djyCBwQq5L7lPvVd3JtGRtLdLhl1agpr
Ycjbe4B+V0Qp7vEl2seDaZqaoaAIuq6mIgKRutXAG+YZl8RXLJ8lukZbZzn5e31Y
2sfJWPjVcTBAeFrwUh0lpSXOWIHP1kGOOzSuNDA32LtAVmnbbdz+Bb9scYvQU6/y
s5vmBrcptbpF7kzye+Kp7xC1dQKdXyaMYbvpKml7a6q9DokfN+4prJXt0ZSBXJ4W
ybAQKG14YRpnOyNfNHEKOT5ycby2S1GMDlpcSkO3oRFBbcN6GG+nBspYMxJQtgVW
b3dtfeoZVn/yToOCJKKyZTR/HJz474dcdRWQ/RVx/I+UDXNzf4G90RTBEQHy2EU+
5UHa/oal+6Obg1AD0KlP8BipTfQemk6hOosxgz/9WmG3hm2j9y9F2kwXas8FBx3C
3E2TKiGdZ7IKvvspNEI1b8flzc7ua26V5A0znbwB/VkrH7bIHz5iYbopER2MXLqH
ljnbCvB8yBwD01eDIr5jiuYGZRfpR21efGe1FAcJHd1WV8tEJYgzOWIlvLdOxoBj
SatijRfcXHIlUOyEJl7FCpswq2ZiZcHXAWjifPYQwDVfHPTH6PuWetJ1e44BEHZC
L31lyKwc5E7X16T/8ZxpJu9VJlvQwacqfQfRYbkuyeKimswgxcHe2Dbyb5I2Jprx
3VnyVV2zJ6o/YOsQSY1EOHisIrTGaQuqizL7ZrWpSLseC20t0+M3NUNcUW3G8E1K
jcOc3/Qm3z1WPQ2T2pQpAkie4mYU50vMW62h/m/eY3RIlYOyVCdTl7pcQhLZbn48
e/V3D6Yz376D7oWp0DLGLRDGQXWqm/1VmAlBO87vPaG2vo02likqeK/KdI+87mXE
lG+Zz2rVKfbe1TcLCGvzn8xNBF4RE4trYN8qKShBs+7Ib54e2F/sJneb/26qhI2r
xe2etbP0nejUyhh99jnsbHhvJ0rHLLSc+zR/RIZAHCbCnQzRFoiCHH5R7nP6psg3
Euieu9nrtZTPYHXLLbOTItfwJlFy7/5s7a8PzDHk6GTOCZtTonDThPkM9oD3cHfo
AwTr2v6yJqgxheX6FzIlSD+iwvkTgy3NlBJgbSwBMRHzvKZz371nGedeTwdAf1BF
VhB2ybrh4Cs9OK3wwuzGbusVW+f3auotfr9GDqYAxV3bgczCMRIyj0yDwRAYiAUF
niTSAt8FGa1Nw4N9XMRr90cvB6BgfqyOLYHBTn0dsVXmAgpnli1VF4vl6hquUvaz
fqBib3sJsuiuz7Wjtskvt2zU69PuPjUJjrNSfpDPB9UoUzxzoMIt5w/SR04W53r5
dxV3BNX4l5Ci5RYmMRRFf7JNuvDgsjTeo/2xbZaQK/FG1nag59oyx4JZZZU/Z+FO
qGjcGqmCNInk4aBTNa1ZOp7cp6vu2P/onJ5rmzlOIWJbZ45B444rfNejcPpcuBW+
t08hOiVSna5wR7q47M9iNxILSNJquzOp4mI51nKW6VdRMClNY+Vl+TRIm5pHpNBT
kqV88oP4mSLaqzsxZI5vcm+PDa2obtMp7ZUabmKGWQ6vI7/Vxms1Ra1VjOKJhEDL
H60oWm0igX8YBMJ8YDr+5/y4p9KhJiGyjqRzAAq3jAS7scty7rrSlpPX1/BVTc63
+uO8mhsEXXqGq0/m485jcyf2vGJMiSN+f7cu+baoHz4swAMFgcxrz54Kt7mFZWGe
LrXwmQw6dVT6COhXVAAT85dzh+fA1WMaAEmuf4d0rTpO32Fxt1qyGBaFD53cgBiR
sgaD7Mu/ulG/5TP/oTBLlzTPR2YONwFF1GD/iqkF9tgnvTTguu7mSGqV0YaxMc/B
rAy2TH6srCI5qeqjmfxhwu5GvrQZezNglGlBptyYZyjUxyHk9SX9hnGSygwnC76v
qq0F0q6DoMit8Dfdch4aWdrZ39H06Nok1wHUqd6gxD8KDTFLhXS4RDzXiuAph2h5
Hyc+P9AHA/1N5p1iNSoBZFwyurgn6WyssL6Swcdq29MzNhlnlWL6MWHOrYI2/GGD
xFEuo+wlWbeFk5Xj9BWoXs51VJZkLMs9YuW6a15YjfpX5hmhTDzOPRgNEJn+D1SD
0RM4dI7cRD9qddT985pKvnc/G+ZP5pwVlb6VYY9ejG2dhdomKxxWLMRtE7K6H4Fh
HK3yeLB6AzuRaSl6fxbgvqMmG4SM4nRnbImIdMqdfNkH58hp1Hvx+Vupp1uyFXKV
GtUNxVqqffEStI0Uhmlw2gUen+Md82a+EEHshz0zWWi+sdfMovlbfmXlk7HKnd83
h+SAnO6CtYph7Y1u7jo0kcKrmjOG2O7pKgcI7htFsy+1b1CwVQnmTdJq3gvu7Paz
SitA4EA8xOpP266Luc3UM2eVZTKOCA7LZEPVs9ppeRo1uGf25fd0IgSPjvCBIo+i
HEEFqInsPsMqHZwt8e/Hj9GoEXiAQ1z0/mphuHxh74o5P/l//zD/rBCH878IWY7Z
rN7GRHkzDP+Fmvk/GdJM1vqQbUMyLvQvDe3ZKWT3KbX5l/tR/P/8f4HuNTGc3I+z
MTqOlSNHGnkCZFzh17PsgIZE6ys0zH7q57UAPyH2cYbErC4qjvJIwq1VJW0L9oie
nYZ42P3dv2AAb25WXLGCOsAByv4sRn23R42qpSVIflufW46VXHRmA239gWdwnmvc
ZWJYcY38ch+Nw+cxySTC4hBXusoIT/JLmpfm1PCFGzZD2gTXoiUj3fLVDddWs51w
/T5PtE3wo5F069iAFId0pPI5345VoXaWmKrN8CrqmEuLTda+MZLOQJkOMuiUJm3Z
lGPDJLgDscx4iUjxgme5LvcgKoffpC05Enr7mlMWlNo/Dzj/9HWhAGkSjV66thrF
AtANR41tnBPCfEnLBBXtZpALBpt49P+r7iXCNyvOyv7atVynn8FP8a5TuIVwbkYo
QjsX7uIyFcKwiJIobkwqtXgjO+XuZtKctB8FWnmWrhBgkPLNvJoIlsLqgMaySqFj
w4tBaRtmEs77YI+do8eDWhXel4aDuzH5qfcbMJfOcvZSfMNIeAHh5HYXu9py2toN
aNGl0kSyoPEnNgDBx1qT1ci00pcv7ehkq7OKtQwVQBFHQ6WTM6REwznR7231rtwO
K7Yex4CHTG95bsgiycDVrfiz6sFduK0iUf3OGBftFx28sTQokVMDSinidu51DClD
RQBj8tzy5NfTwBX/JahbI5XqscX7DDfCSx1gLxQSjeHwNdrCRb1GSszESMbuUqZF
wASvC4I1r0jXCaVGmRQpPtlipzsN6C/4AJkgxkGkEg89hV6qOBvgesttXUc9BISm
DYaN5hAOtnBilHPIMvdmVofB1TFW4Nd6jW47sWwForvCOnu3ctTtGUzwzhV46xfs
U1Q78Rnyn3Mc5z8fh0xfiw8PA6xOJPnxPcvN7xfCPTJe46qCI5LpAWjNwck/sCxL
7noUSMBKzbBYGF6piBJmkbQ09nwbid4AC8C7MBBz+Oa6Bee6hMxih4inXhau3v5c
JvEtahH1qazS2yXqtk5U8ST1eRoXF0utN4xOBn/vw+tCBw1+zpOyaExjIp0K4AQ4
fIuebyy8QoOjp9HwaWSrSeuYmMPyQ6KdFD9JgaQeJ5Bcz0WYkjh7gu5M/U2uKpXK
CeoAJBfD4i4V3PEkvGWtaSsKxuwCqIzD+Ak4YRX9XbOPFH/1Dca/unxe4WVkclIn
t8BR4kWFwidaWtDWTu+VPeUx+IW/cUL4t7z2u5Mf7GmfxLybMOqolwjfCOXufxEw
YOOC5ae0bRd927EQRzXkyF/+LXU/QpIBZFMwm58qFrwUht4OT6l5L9s16fE+5IX7
fi50QbDTstK7FA0yFizrcN1gdMgzNBBSmqJ224qSNgKPXFPJAULA+qmIQnx0Or4/
lpSD9vhBVdrK6BKMeIZAaqKZgIyiwJ27D2awTR3h9Ic7Htc1VCPTp4bSWxn2jj6s
pdVVPY58RWqWB3SxvpYG2aTovvougL1JluN8m4GlNBVOOSmyr6crNzh6BIRmCdpP
hFeerZrRsR0HvZ/45CSjASEk0OyyoF4IRY+DlHEksWPm/eUZ1F0zGzgkb5totn5y
v4f2Z0fveDtI+u3YJWsRH0oaDJQP02WqDze0lfvSBuwxUwf29GubExqWoOEJOvhu
spFwrBMhBk0ejFmIxtKw0OKMMqFVpja6DHiYNL4C+5NQXBmMKM1v9kCECHJJmeRB
utAtU8oWGat5xoxrqzE6ipjZJt0Sgla5qF1OXYqDBvVfDgK8ZvklsOgzx5S08oEu
OCCOdQta9Bo9WOo6KJI5nwgxIEDeR0wzBs9JJc7wuxoG4Dt2hIMuVaSDDUoqgzUS
PJSS7aHB1YZWFSzLG5qCComZF/e5xNtpuaQ/1ghcJ7FyFm1fO6fojszdaS626y42
j6jPQQ1Ux962zpM+URP88ewdRni/I0tR2/4Jq/+MyZHru+9w8P/vTvhyc7lU13NN
C2xg8BN3CA2Nlz0RfSK6dGiTvaix2DjeSjKjjOPXdTVExf88Rj/RYbPpQMT7kX8C
hLXnvi8Pa/6Wa1xjUgNFeoTgzhb4OCfN+aopxPWH43NPV13vZVoKPUYJJHC0qckQ
+CtaHWgOdxrPkh2zQg3uCDhwiDXEJAadKfIvX2Y0Y5OTgHKkatVfBZi+LVni2QaN
qSav7kgVQnyBRnTUU/4gYM8vjDMcmNawpeEos+3/I8QkYUTWnNiZl+meMBFGxMnS
PpAdCkEnEaqeyQK9WovIIrRjFZJoImEt3Kxzakqe+yI/P5mU5SoR3HEjuUYA3WSY
qKuzMztBRLw9oNnkw/3ROHh/qqEHAws4PEY6Gwimxeq8pkO0cTJR4St9T5h7FQ5R
s59vPaeI1oKhBb/V+0RZdTQh83mpw96JtH2IDM/OqrfznT1Ky/LAUaPWXCGKKOQw
1pEcNayU18jrFFwdVMvf2x6TgKA6q6GGLhgA4GNhut+38kTqSkoZ1/beIatjlGd8
fNmtGQxTONReD3V9o/3Cdh93aQitdomeCkGSA3W16JNKJgBM14gwAKIiDE5lb4m9
Qz1hdxByA9bELNPEfQDX0JkL7wpZG5nPt0vgfLZDTAUUVyihXeA2dIxX+k/yHAJX
LhmU3kVMtvVTvzNa1HC8y/5jA6x2mHsARM86tO3w2yJyzbpjXbbQU8F/BNDDaHQH
9hbezCmcCxnFAxw5edgoCn6r89SO1G0iMFSjfiMlovpoly9XRJSp8ila9weCbK37
i3CF7+b8kBnWXA5W3q3RhA7aHMYT8KHK/mWcxwdhT4GAWBfbSTOHBLLV5itTNCQa
qoqpaW5KkYfXTdgZvbA8kgb5vE+Cf59MY5zlLcuQzBmW0GwO9Aee2OHYG/3x7n/3
g1eBeIvwHjrCITh9avwVvam2RbPDnzeBuBSiMd++pmNCxGumQ2DG36auaT7LSJTL
c6wS+wXP3Per8YPl9lkiPj6sAG3MgmI1BRrqvAv9CUBsehn+2ahjY3E1c4SdUY/Z
pKY64cKMSt7fL3c34jiq6Mi/+24fV42mbewV7Nldfqj2BGneBMieFpxeo9PuBa3Y
9CheZ1JNUzNOTrdVHwzSjbdMOuCj7IfZdkwqOWQzMn5SYfXLZ1LhLeYnTNGj/l3L
o2+xEdXPNtEAmSTCyP8FeSUeN0FsECBVS9hrm+ioX7Ktv9y/KAeh0KlDJRPgcFyz
gfDLdYZosEIeK1/kvuvTiAO/C4BupuWQXVAk4o4IYyNzJhhSiLPf+lRNCwV0gc2X
zDvo+pHZuH+UfiBqfnQN44A+RBmi/tmaNRdphuT+MRu3xS5qzieJYEa6Z4tInAWj
vVv99r3W7x7ctAG61Y5cfUE7O2LrPGvtTGDlEWroARhnCLStl+79rCCIK21Tmown
U/9hzc8EuGgjYMp6BSyYsUqU4ecxSc1bJlPs4m7CZs6Zf5uIhG5xs7B96hiEEIzU
r48Vb460RtSiiUeF1VE9Cq3n9NERoLO9O+sgJd9k2fgXn52uJXQ2RbqIHXzX9Hnf
mQiOTclax1PtkT2iRBRVzIUg/LtnVhRSDci3lymSBcG8eLGrMDB46S0HKgglfBTz
otstnBPYXqQRdKqlKGNh/eVhUxhsbXjrZI8JT0h/mIe1LJDO4LnPR0GljGhWY3tr
Ks6JTl8iYIuAbGYagndsCmQOIEuZ+PKmnny1se1usxzqbEZUZR1YpsdkXSs+b99f
XSJWLv26wLswnhz576m04VC1s0dWlp1fZnxrPpltRbun2KgVcrA6C7F820OBkHx/
JSRNJ99wXaIo9gEdSr4CNi6+TAKeppxytZd5uQK/Jr0joJplOJUMZpgwPyOQyG25
CPDaX4zXBSSLoDFzLpOK+BRDHPd94wNFvBoh78Od5DXLGLg3lQc5NvFnlRUA1fNd
QE3E7wplbMNBI2wrrpns3Km78e2cw+UatOFmIK8+fM6LRQ9ZHHEbF7g7SXy/VvNh
v3WgwW5GiPhseutJ9VFnYB+IW8iN+BnC3DPN3HeyysnCCkFmpwk0oG6rfOljWPtd
eU0rVHP9XDNy2gJmkzpJCjCxhcXCsO7qgmmEQZUnRpVVXSTcIVW8FMJcxxp0/Z0A
mjZaPkOSG8pSGartNxKnGv8nSS59//vIZ+y6ZTJReqSUNeua8M96YfNtFu9joQwu
UZOStwUQsxH24L/CC590ITUfRBQ+gXCFRerYacFW4V7ksg2R/Cn4wknbOU0mAysn
qRLOVugh/IiCcXIePIkL5QK4FhOswjx5R5Ik6+CQzHOMZh6SxTljVgSQUEFkLRP5
GidCWu05A8DuFdUFkaFM6yLQ+Vb1gLhNhXH4DyvzE3vQRnKUrfY8j6/CeMQXicnN
EeXecdwZnVXTcyWfzpvHVYXQPGPH1WhyAsH9u0t7V7cFFv/rwLrD7d+rx0TiW0e1
Uj3s2HvWGqaBMguZAVF7LqeHExsMNpbbj1/tbc6OTHOyOO9KlglSBKf8wY6T1pLG
inSI1ip3SjSz7etToPV5Y4oBzm/Kn3bqe8OrnMufE1ItprRwcmKz854QpvVVMDOG
BnFP225AqMvjnQoRbxclMyp2afjlUISJ84UT/3GSu6QlSYm5tdt6tyiWoSfdEYbI
HookPF2z540j0kFzvvBFuPrS9+IUYQ/2mbv2sXuzJq1AEzXIIW4ZDmkQCXtm5EVt
YakNBQNCcQzDVQyHMjxS+diTU30MwapAbUWwFOhcwfkIL4+2X2SQ7w6pPM0eSzbO
LvIOvu915+Ec79qmGdvi/Th1W33imrY0TqdflB8xAKZmVBJ+HNH8YG+m/1p/Z8E8
LTYwt+cfhBy4nhTXa/06sMc1f3uyqANDa55x+RPZyQi/XiCX1DAL4bkSdwV90tUv
oC2iSjE5DkRWKlg7QJbsspJomm7/z9SYlZNZVi3DKtXU9gJnBh/izwYKTVsilTgv
pIHOC8egsdZKoPrYVacrC7ZA4cJ6g2FP3M36W3j11AXU9hAdz5nebf+tswXQIA26
45i7MAqCdlPREkN6jiQ0FD6ZD6G902KjJS6i2VfwuAoLJJbsu5i0GKhe6T9NgQ1S
w7Ig/mc7UJekKrubMHWfRrOvVmWoMewA/Bfn4SKp0aFSDaXyKin4vs5tEEyuhq2t
IvUAfn3Lks5VKCTCXHyVctqXyXudGUZOIpvXBY82zOLs4qufHc7WcGSlRXPcXgaK
JLpUID89rBlKsGvuONwkOPbUEClqHLOvhymd2okHaVh+Lsf27W6k6TV5GMnXTzSU
gvqO2sYMXly1hP270eSxxAeNa2TvXcelJO3gGtP8TtsKbMM12t7AkhZpc+lEdDEp
RmKUU+rYXCP4IBqu/u8SP0ED7fhzh/WYym3JpseoSNo5F1AEDnzdmtfcweJqfTDQ
AxTFmpRjiESIq65J6M2uSWPATGyJPAM3pBYXSeyr0XhSsMRrPEqKzDUWEL/lzJct
Jewo1F7VSEhrsXpQnHmvEDefDS6tBHKD0+kdkY7wjqW2itPKfSqM3WX58rBgmWoA
BEJs1a+Cg7IFR0jcAQ7JQpQbuVnXvgTzImpAq9StjOQmeP+eHpAMcZaQz62FVsl1
17qe+vdF6B7v5fomwwvjTsEH5efQ9CWbYnQLGovEZ+jNjxa0l0iZ8WakJU8x3pQ9
5cy8ejAC7FJte1N/ja6wIynrM2+1QUBehKql6upDkR6ri6p1GF4w/cN4hukFrVqR
jYP8YxL3CfSaVcszloaNjEN0U1D5SuCKj5seQO98Cv61aNTxXlOswmi+BTQjGEEE
Ghhqcvyp3xOffWH2FBpaTQG8SQgJvy9LZCf3k0Ql9pk0LOKZMmYpE7NWTQW++cMi
abi55lm08+jHZLZ8wOKXuJmYuWl3rT2TLlZxTkZ4Sr7qkO6u5yfZGt0/VE4Ms6o+
wfl6ND3Bz0p7yCkYYfISjm6E9PNxL2UEsnYSc3LICDq4NV85+aDvVDLUCwcDMSTv
nZUnt9ldsCbERIqPDvFVpwOioqC5hDaWuxGN5r5Y2LdEOiDuD7570HRPxHHqZ+bW
pAvk8K08GU7uc/MlXm7hmWWcnTAgQ6qln6CFIWN9XGT3vKgzc68lXVW46zrLcXme
GA0sIrKnpogWyieWntZ9F+4lWCLSVWzzd9ifARR5Dpk/a0d+jlL9kg9j+Jg1Iopk
bq+S1ix6Fz7i8Xlbq+RPZasQqjI2ul1fv+5wA+XOMJSpfC4fxxGT42odMwGMi8Iz
ELi3FiFYApCTj7ahs/dde0EpGX4kzcKBQwwkXmE2PLcWsZK7JdpGHZoNlwMMBXuv
/NdmIAAqI/wFQXds2pqWhppJ8nONLwXEhE9eFRaggLWBLwhFeNGH7kcPyps3lTp1
4s9Sm6bCxViwkefByw9ELp6kk1WlcqNyjIVO4xFEIdgotpiS6vzLTojk583w1U89
wZxLXqqTabf1LrnDhKj09E3OuBf+ptUWb+DVgPXk2vTyPs/LCFib0VvkmiLBFtoz
RIQtKnNORlAhltYneXdZ7AsD5Q1cr7dUxE6hJi9gilFEfhlTEWWTE7Hq/Wkd4WFw
FBJ2EEPfIdYwGQVjFxERzEQio3QnNOG1wcV/e74igVFyyPVQdyYjyJxWuB88woAi
RzdTpzExD0Q4iNJliC11N+XztCP4oq2CEY/miasOYUZrDgY9xglY3MJFyFZDIZoU
qtVoysyXOFMjoPaQjLaHbzFT1U+foGpoxqLF8R99Ui3+aKl3uzW7rx0PxZJgEkKa
avlRDJ5tTjKQUx4rObSHI7lJMzKbXNtAxYzP4deQuLEYYsc0aK5Ndzz6rmxh4WLE
hIxOnuzzLxB46+FyYexQBgOC4oESQqhv/+ilE7tlMaseT6KlsCoFDcMtkZEAs0mA
9lEsO2PsUmSRiV7CslrjedhOm4yyLgsvxymjnIiQuXE7aQMMbgmD1NphadC1K0a9
D+S0zU8LSat5IYT6yxiJer+Ky3WonXiEiuO37EyQLD3UtwEHeUwPcj5gYFIrfq8n
92RIllQnS/RCfkUU7jQEXLnXDFAHohwCo68rnqSdkxZzErhNqZxgaIJlqdjaJAhH
gKdQjKnT20GFrEMX7SvfPG/Fh++PRN2CHpWWDsEegO8Q3jnRlnJW3b1ZcXBzQqLf
vyONwzS8d00+YBFBOwIxQv8VV5/ooxtfv8yMBI5wg53qOSHohPc8lKervZZzB8cM
lSBMEpR3yo/AOOjuHM4tFoO2+Ot2IuHOQ6dC/O/K0wTd+yxAAsZ/2p0yPaRecEbd
ymPO/ZEQxFvCpMtvhZ5/50QDCCT612XdgtGjfMdcpUFqFAmGsw1oWoj3Y15edYOz
eA4o2oUYSfK3U4N8t9aJOZJA6KP0NkoFWrxyVnggquHQhwZgMXJvnMKSJq4DAimp
9f+UUlZe4Odn2orEVhNldcCn4p4Tzvq+hMPZ8MqF8pKfZNhqE66PPCpOH/aZihFF
SCtxssdiYwKl98wpUW476hy8PIxvBbQsBvQB83dUiCu2kQkJzAZhkzIK9YzuUPvw
ogEA8lDdsR4RiJQnExYyTG3vfIAdnKZhEYkmLco0el9cJ1WPf2oPiD+CdinMlVU4
VvMzGFJKhjKb21N40UIhSQZ7A/PMB/M4EaQaKOyZeGG5EjgntxFrZO9alb/oU6wP
X1r3MgkHLSP6CrTnfuSRsaeAPKtKFdNpJuj6HSrl7uSNZBpaC/PBjZez2B9zc4OK
AZ8SS2jbHflZGVZFxOH2dNGM4PzvRmYQXxsCYxI7wiskhxT22yveBkbjna7Y5oox
flj2HAO4a55+iTphoamt9hx8Qp5yQNYiGdf/iqesdmbKkRYgEnlcd+o5jp4XbTdg
sM6KcbdVplaxjn1+cdgQlf7Rp4HN4AzYXBz+8cQRkMxPc2vsT6gI6++x14rzvP78
WIq4/PTiZLOpu+itt4TR0AUIFQMXtuSw3UJzIYtigMB8mGMSdmbvJDn/uV9nqdHg
YbsF2zggvrOJaxUYe9tWOPvxoYD8OWc4o7/DQMA2ADN7AqPBKjJUPnmtwquKc6js
CjN1AOwq14r8dswYStx71ZNsH9nlbthh1E/+LPVtNTwXanI8KfJX/QzgiMQ+g8Ox
FssJx16zsmxzZO3FL+qvi9FE6KFVI5hmiNQpn1pIZfZb66fQWcqWkzCBRLX6MgcC
RrH1dt0v+axrf3SGLdGiNy/H+K48TQpK4My94FE56kNFFy8o7lqPEfww+lfppwxa
NF5KQHvIlx2CCWnbXrkmFz7MDBk1/ED9JYgdTyV4XoRZ+lTm8ZnvivrEnwtguXWw
P9WKtbFEJmXj5HGDVEks9TQCHS9An6dA5a4eDgZXyPU/GxD0awPXsoq4vp1+TcCQ
eigt9mZ7GxPYUeMkR0Yw7G5nYuOAe/ZUGYWf1wFAhJ7iDbCHR5JyCQULf9siEBMM
aVc8iMLqt92DSyruFgEgOvn57kyk3xwY+IfwbQmdmsRbst2CQMkLLEwFLP3plpcM
cRHgwFESGJgVJo1f3q4l4UiFi/4D0SM/ukmw89bzgWfSIKcUbJLcuc4z+rc0U6b8
VT+m+tPhNFqcYyxhdrbgRhyB1NCl0s8MJOTac+I8NdHTTEzzv3K3AtyIr6Zffn3+
R8jVOsZjqmumwIfFiqCwjRfBaRTKC7TT6bwiFCYwvRwRSN/mvejOfAxWceVOs+Hv
O/qXnUmrMazMD8OtpDbaobTsW3+RVRt7U6Dg3UzGcBvteP8Un2pqVjvD2H4luqAQ
yORk4uQyKtH9tJvr9lguOrqROMutgGfKXuFJqpmsYzYw7FVcXL7xNarzW4ZkDmtS
4lsUjFRieSe8Ls01kJfEIZJRL35YFCOm6fDEs4zSNayuP1wfzrBIQpKtX8q1dh00
E0ZAyD6mvlBbVVBL2k6XXikv5HyWxDJbfYsV8oXF7d0TMmsUfgJ41inlUw2QY0hI
TAPmjIcbYCvPXRaIeUtHc1dLHSmxw/eSKdO564+z/kSxN0dM0Gj85sy1IkfYWZiZ
zhsNRal7H7+nAwmF6+Yh4qJrbI9ZCa1PCpXTRe+RD/ZMDY+UDxnKttW+89ukfuOT
M+A3LrECP3cipYM8VwXrm9V9OQsEUNMhH1GdsxGGq1m/VC63NVXakPjj4DKXthfE
9weUZaO5jGiX8+smoyF9aH7KV28rWVUN8no7mqos8mLwB0cT0ctjnulgPpDPWrVK
zV+sECLgANZ31I8f2mfMrkYoPQkE4Yuca8kIYhYyV0841TQqTkeKbu/ycchtI/CE
SD5Ov+ke6op693GYQQ+0jrn1M5jZvd/Ta7ZNWsKSaJbdc/KiV9QTv/EAIPV79ih0
rCAYxcxn+uu/bBeC4fo2I+SFa3aQ5EE4gQbbxKPDKmPHRwgrVSpipt6Ti7XFxJax
5sKkV1WnVGA3ULBQLXNMMARTwIvdpmLjwPXBDHq4qx0hPHec4mhqlvylHorSnxd/
JwgZoZFFQfVv+G3EdpkxEGj04wUJQAawUcYiw3RSw6uy7IOYBC4RC2kYbOgaCwxA
qOG3Dv54AeVeeaQLI9gqoQz4IZMFdU3IwEvomT46rUOhd6XbtQKhG1WD5l+QrxpR
isQAjjWoliDFIAT7kXWhEFbBNkaciUd/SprPdDebEymk4jYy1hE3zu2VzTPBIyvi
g0RzLEiT31PxPJZh0bOaKdKa23FZSzNp97nuyYWda4GgelQFBP+vvFVHAhLVj03l
0+9a25PNb58w8SCpuHOOfwyJndutHjHh5d4OrMifx1OGbPvUsfBEw/xuwETI8xeb
VC5SnEkmAOFZ5Fu3MfSk9rtsM5P9QB3h7uFLxwW3cmkZfvT5LaD8fHLL40d7a4Gy
3brdfx3EMfp70rxTh/CdNA8N72VZ3QEoxxRimpoJ+P149PLE8mkqchIs2Id0sbrH
RvUV/kshN1ROywHb3I+rxnWX8ZzHkHzFICWZ/x3fqj1OCjLx6ztkp/dmBLwzxtPe
TKbmuvu0ABfHsUnxwrr4axpwa5MeygXEvLGmqWC+MUhhL2QgVR0iydJVSO9jqB4F
0CH1NkPNUYqx4yChWE+5i1Y56sm/KTelzpXQmgVpAHN7eawYERNr8QRkp0mg+FAo
J/YGEGbjgGSHuobifOiYuRcDfMwzn0wb2c05YnuRL34DDzk8RYf+lpYsMUFvkQhU
SoY81jx2fr3+9aOSjJCU+xJxuxrx59WijGCFQSLREj1fiCk19PKK9uragqFzO2uO
3H2WXaKxIetjldAYSsNzoxKJZVlN69+L79/QVEtdYgyTqOrXj3kJpUvbvLAQwniz
tLQJPxOG9EhyZuC3L1wrfYLVTY6QIclxo86hlQdQnigk7lDm/RpA/hghPuiWXNAC
GIjdGNl4WLDmjjhx1dsYpWEDq3Hc9/fkKTOkVr7XZp3I5NOcGZTxy4QXqg4xTH6i
I/Ke9PzZYAsp3/XTENZ5J6LTUh8lRt0U71aywbLKhYnayiEGHcpPEeXpu/rfRxDK
qZsB8OWJDfcuOprlK0yBNIwyWbt4KpAQ/QaoM+vCH5J96jewSkKgi2PLh66bHu5u
vOAY/bBHhQauwVBJYLzsM84Vy+mZAHb9j4pAxHRWZTRMlpPpxN/Ex/8bCnm7UR3p
ZMF3ndtTZpXtZsbVEkhl/2tRpdq/PtkDTTh2PIeYuJ1jNRXlU2Mf2ozNOqndZKUB
NIBhVT9ikq9DekkOY/iPLREep5g99MeRNNdKLG69nr80ZH93HatCPrp2Y8AdFOaD
UZvX7F/0D/aQQRyg3ZIGb0p7rNDvvPzX66OQHxyhMFtL5vfhH3fkFnhWCAoDL1NN
RmXPeanktGGP2w62C+7tB97VTkVbcVeAq79yNQjq4/xUb/3KZjeQYgkkN7qFupZi
aXd1jliFwuliybVm4gmel3JDBm8BvwesqCj9M70ljXmfPlpdzk1Nl2Kess4pMJDK
m5c8hj/sMGHH6uCyNE8F6OtRQtEHz6DJodX/7AuN/HsBreA9Tmhk9ZNLMU+Epot+
piR1CHB2wxse1Mt4szFRkNIkBXnR77D+XR/gczrH7h1/JEodRXAGooZX8mwmEO8i
HL18Vt2sIVnI9Zq4D4Icac4sZbnBMReNNE1YbE6c+O0uz2PFrth9ZXsOuiFOv1BE
DqWEmAex0Go8bp4t0HTtQrqzNHdg/gBUVzMlSGZ1OH8rI7UILepJelO+3cIfAMm7
U3ZK5FGFt69jduD11R1Ak2I0FNmgymxDgjm++yN+MmJUM38HH5O4kylvdh2oXJpV
FadrGnR2X+/lHXiXz16rsNxqE8VDbHrFIILqY2XeOLO5T5KTnTE31oA0kQVhi5WS
jSRpGoeGp/ZklAH8NARYSGCeIoiVjkrit43L9OkZnQZILXyYXllBe3GwGRUCrJmQ
DkJWMpY3g4FDu8Mpr6Jxr9yl+YefaUlWO6Vqfj6719JqBUlePtQHf1LtIqPZkrPi
wzF7rebcHFyR/z9PmQAcx8qEiWHH5Io4wF/EP+Gf3Z3guHfWUM5LRkc7Mi2kIZ6p
kgydzoy04cVVVcGTWCP/1fawKlDh4k8L7pPI93vAGWgBWXqba1zxzUwZQ52OzO1O
Ij4HfuSh2sidY29aDlJzOkJPOHPSIkXGilBZomqtkVgxYMDkMFNxAqGhRuTXcsa3
WH+9LNSSWHWCqoy4VQON2eJvxlw4+O+h8rruVTKLOgRwrqcY60Va1aSG1chqDHk9
NjHzeDR+qLNYjhtG6cQwgUIlMUM8AoX7lRcKj56/cvyqabCdoqbfDsTa11MrHAgm
rwgXo66zUivVZhrfz74qbewOw99NtixzEyLYWXdMCTXaYFSIGhtW1vwWFerY2HEP
wIaQRyihy5zopEN9kj8VVrTsA9sRrtPwebNKfdgPKLYQ38fsPwMaCMi/ldURrVGL
4ldgLi5NASeyWsNH3srgp8eGV89KHHdi8jWpFhdxKcz++AL6oBYqsrUiNOLCMsUM
LUrPIu8xd/Z0db/OpItTMWKMQq0XfLDq0daE3h5vlPRzhN1wOjXHbQNNaReU8JjY
HYBT3jsRdYji4PW3P5vpZCi8Bih2zVQtDYmt6ypZtb8yxqq8XPRighlUc3MlFks2
BSLUslP65et3LN5p/ftqtmF5HxWEYHNV7GjjnZrHVa9FQQR1fCs5oLt+HaVNo3Wa
zUp49cMjeeSJMi9x3waxcmf+rINmLz+qSvqPeYSByYRvX+80ywkVSWTIe25gK1ft
anCXLJZOF7ZKUlZId/bJh+s2+S3BEqkeZ20mwZmdq30oIrufWW7Nm7EqZm3ibs4u
1H4QesDwwKKf/f+k0usO1ITd7U8+AxrJMugSZUnmrL7fXviXbcT9Jm/MUTii/XUt
JYGh8r4tDoYdHHOkR1mYFqee05x89kMeCJS8AlHN45jFcIIa4PLjk/1F6zKn8P4c
s2sXrJ7GI1vzE+N3SsVtmd0H1jJ/lEqffoDwZg4OhyJLUvfS4rbN9GPc5uQbILwt
IZs/6YlSOph/GrKXQMn6oEyKC0br38wH3Fa6o+jzuV+JXtczJ8pxq685INxc+CfH
bvBcjLjR/obJG29RE9edcBURcYBCzxXAxTVmoe23wt7fAHL03gWPjPe0SO7FGhqG
faclbfq8UgztkZ375bYeuRG8G4WrMV7wXRWVqBT+sMcZJT1RB7cAJ54/anW3ymHp
Q1NZEmOKRpA05TMqXzIx5TENRf9gNcJGEldVCTVLizZ2pyPHYfdarfmf6QDtQPWf
4brt6NrBQ+xyrjO6JASLlWeSVlIwgBztv8e6C4Y9vikKLndDiPj7VJ3nuT5hqv2M
lVU4ZhLiG7UO3afXdOqUFbGZDCM6cXkahFWa/HXtSap6acSnSlB2khkdqPjK/vZ3
U1zD04VlQK2ih7UQ8C5H3rvFjBGkw7ZZPB/tOBw6oPcoY+suAVv14rOpZlkaOQKw
88Ff6gkxmj9IlH+O0jO7tEd1olr8E42Oc4QWJ4z0QmdQPrKJ2zFz62KL8DXag7u5
1+AxWB7PjxYiq+EDckn0gkPwg2byIfvDrdj1Z5uK8V9USwEd7FjUlZx6uoSeOoxR
x00r61RZuGrfGXtEBPe5JaDeh1RDvxbe1jcglCZOzKMM1EESexWJDlI/v4TZVa+9
PEPc6x8Z69hCc8W3DK+kgoMMdmQ9kVzLQqbJRSKOQBYS+0ae8z8VT7R+lHQPTHor
glOMomPcRtgHzE1tDQJ3Fi1ZrhLNmlmGe4pMDwZ8esw2IgcMbTyLGMimRIlKow7a
faIiyQZURDDPSGIKVcEPAwXQpsTFZQCN/PbWcE9VlUjVYdBSsX9Syq2aouM3YDdq
fH1LKq0KBgjr22WBVVkVXrHOUWcUM4FRP25NxhQor/Rih83JCDcOo66qe3tI0/Le
RQ/edtwyMSQ4VDzTIg2JV0GWHwBK5sYWZnjtDllTDUMKbo7IIFxScT0JZL4OA55f
4pxtyJOJk+kqFQa6U/E1M519MgvX7+HZJJoUCzSRXs1spwcN8gIspsOUDjFayKk7
ZSPWYGTpZR0kGX7dPdTnuP2fcVYEWjOilCSk02VENw4nTdZxSpN3W7t+1CbtVIZS
1/vnie1G9EWWKO9NrlM2igl3orT/7FTYJDmyzSxEyBHfuOlokOybDRwYz5WbMwf4
pTecrMACX/UB1+Hs8YpFC44RFrYUcMY+m4ey1yM41EXgm88nV7EzK9xu5BcU94P1
kuOLZ/XF4tGZ/ODKupwxAaXx6THXhoJ/tdF19L/8HiVVz0SbRVEs0fly/UlxpNuQ
12s+CTJj4vqANbdQ1p3B2Tn+o5IdGLZoHZNqEcc7U63/+gCwv9CstwsIRkA5CEk7
F0zQwLCxbyYGV/gnw5VYpdJahmHMLmDof4PCTEtFiTqEh8vBKGc+q415cw1jz6r7
Bg0pKtKJ1fvD0VKFH1zmoRGCVYTxlKahQwqfDRfGtkw8NXg1ntsDdHd5UPrD0fqC
v/DXJ1dteE8Hw1VVB2VSao/rBnrZFisbJov1z3+qui6JuGS8Ufd6vSTGempTCw8/
Cim1m5hy00acCSNl4T0sdzd2U6tYQ1aWKx3eZG8yFxkD87t0h004jwjW/8BBG4Us
CLOet/Wba3PDI4LOzLhoFaiklX1xLkpMjh6ejMgPXA75JFlpHOJ/cwN4ei4DYeh8
aRBVYCuc5g2UgDxiE8v/3+5otQ3RcI0z0tPQ0rNe0cO733tEtoTA0koGD1zp7NFO
y7tnnanBJ5zQQBgScIje/y4a5bfBPrwI0pYsifyNyQAlMQJtDxiA8R+bgNPvqG9G
7x96M1Ws90ibfAO0MlwkcpQ14HApWueoToGlmopYFEXQvg9tqNtWPW0/iC96MmEG
Ob2cTeE6xrh0px5AfILhn28qn0RI3hETZjK7gsLVbEI9vgCUf0jNpwlYpv7moFFY
8abO3FeshP9oxX/feua5IkATJw5PIKvDnX3+Mk1rFyIHMT6pAex0iW9eFEHVluCw
vIK89QHITPy0qnp4DDS4PPfHbthwha7wgHIJ8tqPkjHGbbfX+nJdJuypWkoXxgUZ
qbC4v2eDfvaJy5rSkS0IKy5qhWyv71ymlzoybDg+Nt2L9dFSinf3nczOiOVxokRf
TEraAf4vsBrkoem+i1K6k/OmSZlBjor/3sEzIoMmS3ymqfYuK6ehzTM0POu6vCB/
uDpKc3L5CtylbGXshiOiuasCvp87rgUJwhUYsDBSilKJ1T/tJhTVlNTsW0mxF5Ik
1f4hF93+8y9xpIdaDFgpgXvK6ul2o/whDLVKu9l9vnnLv/ZBMJlC69Ycbzkg/tZz
tc5NyQtn8ccKI4Rb6qT08V7Fc20GCgiS1rZ7HUFWnvaUMztiYskPMZnLr7pegP2Q
b0wQJQjCgf35voi45oIaHtgbqhP5VTm0Y2oHo1ihDkkXcSd90Ys2qh3bNusp3g6i
M+7/+3R+P4UqS/V7j7wSh1adyTZ1zZahCDx0nX0olfTRg28d0hnZZ8/9m6k9O/7f
kdOQEgFteR3KGBpJMdaeKrXFhkx5pemgjWqC/fxYN2uQuyivznhBE+HeZkRzBS0m
8pOthDKGS8ExE++MBLFrcXqYaXIB3ZaCG4mVuKkwemjTDU9vGkOHcVjajk+UCRtI
uEs8oOPx05GDxZG7c64E1RqSvWFovFv1R1/iPby59RDIcPcDVBgMoOM6iJBxFdmQ
YMOS+jzXGp+AgKIKbftihYcIfoLDS19MzRXYX7OnKhfoGR7K+zj+oZB6lmbJO32O
XeQ6h/YT48CqslGrJ4/wRmu+vDTEDWrD94Xf5sY05kh4a/pgTLwDNL2QTso0NTLw
cyRY0+Hj5OlcZ9sboSvia7lMJoB9zmsD8fwzeegx6D8GoYWqFwis/Bvkp3OzE4Cn
d/gNt0KOcmeYsVN/7PxIfqAhQVWfs7Dhgx4IlA1kc1hoH0qZCa6t4FGnG6URA2Rz
L6q63W5/UpFjfi+/7ipJMhxY/tGFqr8Kv4Yza1ocR4mQWud5UlXur/JN7fxoc0tA
HwK8ZwqetukafGHWCokSkJdoRL22I57O4F4z865B4tGfk7LVqGlVcKxeNY6S2zuc
bblgo2jeZItux8Py+9npvfOVEeUx7QKPdh4DWie/cjIDHhWwwSkpJ49jimBp5acU
PFC425AhYuTKr5NOhiPiDDRrxbjKZ0C62pWkif8blWASkfA8JQDBqyTVB8T6PlDk
4RR91sXn0d/w9qlxQuDke8x4vvC09lF+Imf3vXA/NLOrOH0z/AgTRHqD69dlauxq
cpotU5eVaNVOC+bI6w06CQof4PaE4r4SNwkwczrpvts1iJ2RaoNr6Li5DoqhBWSY
AlpTX+VS9zBMkmgBNHv8WS60MRwngKqwLoS5JHbRqDlmXZEvfc/mHZcQBYvpx4U8
cDakegvpT7CdxXlp4RpqpDVYdqLXpFpUAik0lvakDjeC4US6IyAHWQY5QeAyJKmB
6DQn8II0xi7LrIADj6zdL1Vss3jzpf6nU/LsaB1vtHTgJytIdar0cHQET3ZkEo/A
3KZDhk27wnO7khEyxeI5oVVOKVI2DA1ffmQkkJ8zML9JP37DOHIvlXEjTxQmz9I3
iGbPE+EOLysdppRXxdkH+Opcb4qKZBTNdL/4pjJHJoMxxL1brj6E4yrhxHrTIjCa
MpOqKUX7S70gz15j+RXbMmo02TJ4FNgqM8GDoURGhjxbvDLhi4c2cjgNKmj73Tkc
pu4M+wPQoa1X0UsI/uchWe2c7KNI+pEN2tw+Dy4nW+UzGdaqv+yndBg3sKpPtn+L
kwgF2Gi5TlrEAQjELs5CD4Ll25Msws2XP6siFFxODAqOSGB/3fo69KtjfbFodeWo
pFBiSCeHeJbkBJe1VLGr+1GB+3sCY/od60ASN08zjaXzS/QIodCtM4uwB1x+py5w
2Bcs5wVtSfw0JXlQYZPjTZZOMgRraaiK+B7RPEg2YaV01kl3VIgur9I74+L6jf0o
jyU0a9vT90Ek+2FQL4+Fqv9DO8+9rUyZsIbWDs+rUsO0aMDeBstVzG18aUhfWXkQ
eZAtZ+pnuPNsEl5LKCUd3E/Q8FyDT57IpNWDAgZpEOGGHnRfBET3n6FPUROa7FMG
KVNpgIBnkilYNeyzwTwDu53uHMpD41ZtFnGQujmsEFyhP9DURnZJGjKxQPMozVJW
Jfkj0qL1YitW1SFA01+ZJc83lVVsF8QFnOxefSY5wvYWrTOus0qez5hLTeD9erQg
mG3WHN+ROJeDpbWkN1mu9Gd05xc9fd+EOQf5UIDmgeaxE/WPxRXWwtLC0iWNy9Y7
6fRZPw6sjWzP1NX71xq4/cPKT6yUlur9bARDC4idON6Xs+apxVZEswtn+BbJWIIr
zjFcydwrilZIftRZYPOE+1uTLL38XCiOH4VAmydSjSxhrR2/ameIGm89AWt8uNAB
oYBzUnnXC0ovt8nBdZ9y3fdbX82zt6KNE2/n0S2tRfcgr9gpKsaCPpAI+XFSMltc
JxTYajjtvOp8/mTgV0a4cl3TGMQtuusdRhLE79VTrUj62NK5/hvdX1exPE6EnUqG
UfGBiihQnl/Z1jLP9vxP94BKVFBy5jttS0Tp/4dK5irG8wXhnqP6e1BDZfBsZ07c
wxDaHFCJGywwOsThhUPIaTiLdlhgQ+I6nkaf+Z2Bw0l+PBs+Apthgj8Y3iCxilpN
22RNCBf0r/8LMPe0A0GSLr9p0hkByAGnFlD8ll+cS4+snnJcpmVQTXIstrwKXdb2
BE1KR7+6Xhiy0H5jp/sPJ8OT4NfK4JCgAlKRdTvp0QeL961wqgMDhNYmq8SD2Cbo
OvhG2SCcqmTpiPOSB4g1anzS6J7mKE5T5X+CuzXWPTbjnkenc8++yAm7hAVi2Eja
ksuqy9hCJzGz1G7d2D5eriWKr7/LZoa8EhcP3NDvQEaretBY0dyE+imsblpXHJd+
M9IFCZr8Z3ml1w+o5ZJkMEuBIywBxBgMbc4NWWXnoSs6bT3ZWJGmrzVgmh5LaRJD
i9RtN4m1LyW8NFvcvu5Vt8rIlAq3Newae0UokgY1s0bYJKyOg1iOwpa8hssSVLz8
sdZPBnWRSzpHa+CxTJcIA0mvEMaiehAtzFMeKVb4DsCI20EvuVRjVBozjVGLqVU3
+wzkT5aFxpu79s3lLWMqL7bn4XNK6oyBN1dehmmci5OpAZrBVK8EEiK3GnwxmWdV
2fQKXOdrMCePjg8wZ6L0MvKXPTljheQ03EaJT+AppNedpncGgYGQatl8J28QrDtn
MPMBrXktdrj5lw+gzi28sLGsaJR+0GleNWaaZfeWoqQ9TEvH+feCzb2KI0lFYw6v
wu7YhqInTTb87rvzbKLeP7pv+OmvABUcp5eTHthg5qJa69EJIqfEhVrMMaCBZt2b
DZ6pSDxkjL5BBhtSI/Va/OPdmfso8WswE6ZplZGjOl8Y+p0+fD4KEjhIOvqBB1xQ
9mpP687z1Yruehhm7IBV5xhg8q3UC3DciFn8IF4jFbM=
`protect end_protected