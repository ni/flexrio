`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 5040 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
KKcya8NExyVaoCvctjWPKTsPXcyaCEs1iPzGnPO3NyiERDjwV5SmTV8rqM5k93pj
o8yQR00tVSEHrUsHrdKPFyoCeSArSYQlAqmbppj12hUX6PzUiNsVgs+14MP4cHzd
LFftjdd0sG4jmtaNhlQASbL3nP26kalAJe/C/kBcsK+2OMn57jsdaMB6JE5gvjY2
e3QUkjFufzfq1pLCoi2ksuenkF9hV+JDxo3e7lnc7I9nViwZUUkzSJOqJfrBGN+X
HJ6J+2RqiTn02zy//CUqknYejvUz8ldClfkxMoFcY4CWUtf/Ybr3KO6fgrpWxva+
RgAd+d1QwYsIEUcyCKccvKqJKDNOLQBSDH57/po2M08j7wMV2x+yOE5ZzBy6b60M
HsanjSsGJaSJKbxHJH+M67UHc3HEAzGDsrHPlNNSWADgeTfqvdF3tsU6Lw/7C/Ih
e97fymF50sdqvM4pyjogCh7zpVJ3+t6ckMIQVNaiHUvRwqvBFwZjKRPb7QzO4nN/
Sc1kbk2XEw+K/iIGPsdm8fvhkJPcxVG7cV/rxJwG0xfBOcU6Y0rQLv0qfCBe1oEN
vYEDU0Oz9gUHgTWS0g7NVu8wJuEoVHJUw5VARbFLlq+BXhpBnsxTf7DIj9RE9Dxy
JOV6VRrr0J4eYblZmenbMAU9KjSwNoVg8QXuhFCeyImInf+U/BQKHiWLGXJFC0+o
j9m1NUrQiLHtFF9v9dunwYaU3E+P5XVnQuy1UNpEKYKs6ZF6bswfJiso4gOqU42k
v/xfMw8gLyu2+Q1KbcustwYgdMFuBYSLyMcz48cR34zGTqMGYeIJg+d2ZsIMNn6w
8FwRua2MuYK2Le2eG2olIODoDvmBdL4ao1nK8kp+brCQPJWdqDVZcSV1RZ/+j+PZ
zczBGcyuHYL+SQtnq7VmYhCnOvbiFAhynEDScMG2AK5v5cGZS+Q044elDgV3EtI8
t6ALvRY4eyZ/VZ0FXYNyuCTb0aSx4fXj+zzYt6eZ5gbOG6TRp2gMsZUEbj1DDZDF
e9zvKS7/niPhXN0yAgYs/j5QbX22D7FXtZeQweyswn29qnEe5u49JIIXn5YpoZnP
scjp8Rh/ZRyaGz8jcVjkOm40xomEqOyy5gLLQlLNrJbrwVzNUFqcZNSMhGGbAqqQ
z6PZ5zazUBMjLiDK3/xBoWZTNrxhW4pzxG+39bMxQHvFTteoovkZ1Dh6W6Uc5S/P
FLznUmuXxkxJBo+yZDy/QNMi7O9LanFQ7SIXXRb46b7UCnEV9I1zs02gznOhb5uk
jSXwVpBqlFrG11hfwH+xez8VXWA+3S9VUOFmSwcuOegI3H+A2FmwVONCInWrANsM
Z80p4iKcA4zM1jZdNo5x+VDirQ57wXmnPeernwkoewkoFwff4YzVdYeGyDHc0PsZ
Uje2bSXpAA0BI2wjUIv3AExk/sLuNm62texRVwbhGdObKXT7DZ1kZB7egaitpFse
ghZGbSLgyrchH/lCD8R6xiiJEpMwZLkxOMsVZYUAB5uO6NfUqzSiIaB/sIjois34
WjwWocmcfldhuAJ1WEACxQ6noFKAy+EMFFHx+8Vdpcj8wgzVxwOKGTdz0XLjKCyd
UIOMzniTHqhd1C4RLG2K/qEC2yQSm72P/nVmuViDZavlHcZjmLG8RD4ydXeliQ7G
FfZsax1MeeiRPK4QNB8aDU4DgkB8e8hLqcCR5EQ5iP3QduHbcREO0yTQS76FJr0Y
0GaMtlceASJbAiZFgjxlslmpueRb+HixrTUhCt43yFOei5tM8E2LMHc9kv0cKemf
CuhoZXWI/gR/JK+MtSApnCu6hYecuVqHEZ3j5OmQokxbg5gWlRys/f7nTNQKgJTQ
S54QtcqlAHnYmCoImq/BaUrbXo2MkGcYZuG/Gg7UeBjmUw7KQt5yAxoQZUrX1hwx
rlQFXuM5TZFYMeaAbUwTnENbxat+Fn8c5nw/1Jxx06R/4ibFIBMJlNYp1lQcdylL
lWkaNEYVbLTKJhB+faTR+sHQ7YuZzdp/yC235sMeXDFdcd47mop38FPqR/i3wwsn
LAUNdXnR2Yb47Z+F3WJYnH+Bt0JHBBXqskfbS5kXJq7exxO3qw1dF5YI5ecbw35k
aDgRpxYZ3CA2K1qdAS6OLznaV8QB2FcH19QCLUdZxneUBPm4k+J3ZOnu9TPGTn44
cv5m6ZMNXLPvsNBZXiY7cs0FV+yY9mRfcxuKBkrhCoeYjM6b7NdNCIRjk2Vd9BKv
hwP4/3g7BhnFAob3lgZeFia+T4Q7U9CAcJuCHUd/XEl4nMu26alqXsFFhmBtVcHy
q5XYlusMlHMlpCGLgZAV6Te9uSfMlUGLvPSAEcDFsQh2CvSler0GQSfjhi7XkkJS
AErZzhBD3aa+fElqi48693i1bvtPhxAmLa1E+gF3PAlUfVR2g9gmzAwYkUeL9DQu
VFHQh0JzjnwK/HSRZAgsXPaKXAGR3aJ3pLNJYFcNWFCorYLucbdz1mJvAANiPlxf
Dv2EO0Jiti3tM1WYYLp6JpMSCRDaH9eJ/O0vR56V3WCgM/8ChGzH78ab4xG46/w2
xb4tRBb76e1WG+KeL9EjcC4lCdhreoj/kbPhSsCDmPqLLucxV/stv66rEsvQDJos
u/Z+UrzkYJ3P7YmrV/1OH1Dv755oDQSBTck/QiZOdet7dPDfTvKKNQn2i4TWoQ3g
aOtWCiX3rWjr8hOF0E9sPsXmSH+ECbkOY7srfpGh5EpP7E0sIO8ZY7RE1rLpZJ3J
+1ficB2hU8dtZM/l9o8X5uZVIO+RWmNo98UDvJ5R75I09WlqKT/gHRqhkZrzZuTr
my3oSw0aubwbpMagy5L0B7fvMI2WEdOjVKx5A2y/uaVym6uCHdZmbpihH+WaL+W7
JKCUeVfDT8pP+HYApwo43lFk4M+lvUb/byN9dlQLjB/rToC4KBA/Ezp9R3m1zqv2
XuO+VlmSHR2b20LuLSHI/mgNt2vOVWFGJ9QPMPhDk2rxRb4y1bH74fVT1sY6siHK
1zb/JMEz6PbgcwEgGbjxQS7uSAfwUiHsXFgk2ZkWr39iUYq2edMg1INik/G3AQO/
8SLOgKFYbyYNWuvvej8fzYsXNBM7vmVRkD3DHR01sU4zFmKu9NWayyHeJD/JG26g
37IYA9DeOwaqVf2F/sAioIzxv9HKNethI0EG11O8uJcNrM2fcO+y7+Kv8bZZR4TC
DKgYNdIqJsTjJUBn8pB/AhW2U5cPNKsMca4CAyRYGXLVa+M5b9GTtUkItpYgqvOd
hKaQLSCMMf4xTsqJOu0WIQK+wkRCJdue4Bn1PWrRYUKiltdKxlSQdMvTDdhJFQxl
Ec+L/boDxuVdK/ap8nAkqTQgsFo55Xhb3Pwa6qqcnJ2YNa1SdZDgMRt4NkkK0flF
/93PL/E5OJYTlw44Tiy0pf+SGAjucURv3ZN3px7ZsEjQ4rlXWNioL1tnkmUbtvOD
XJhLLu/el0+N6Ef9YEXBMPWNY1UiPk/tI8K2G0G8SS41XO2fgrU9R3bGo3P57pvN
OCFJX/yBzle7/SfPFLVQHq++qnrTt108D2SMzfipCRHQG9Bt+cBCLBF3jMbMrtDw
2SUQyP6vpNvtV553V+tdcJbXDnFZN6e3P0PH1jm8WjA6tt7mBTjk1hl5emWGW5zx
DtBC3WxUo7ACGgI6dehnImfUBQsMo1t+dbGQltYjOfL2IfidxFFWgEJFCofBoSqB
CXFeTvsYke7o9TxE8ZKiqUp3TCn73+irLIXTP5oGpHVaKW4tkWg5fteGdyBl0slk
csfU4O+Z1+bsPUgSIHLZETn1lYVwQJjk8cggh2zOs5We3p/4dghvTDgX36/njAJ7
zonUf9iLp2EF2dIbIj4QBtk/5SaHTDmqZhClGZzKx6hDp94ioej7VvUUtNYAvVvl
G/Sgwp8547sEDBB5R2jzdiTvJriX0s7jwKKTnc+OMYpoLjk25Vg64V2LMkPN7qRi
xW2uWF7TwhKwbaYYIRFVyCxGs86Z0ZaGFsmLvBYB3Y2w+Tgu95SsxJ6xBbDT9kc9
+f9nOWihmvt6+yUJzNQZs1+V82hiX9lcmDI5T7Qi962GJJyERPvm5Nog6dqvqJqi
qebsqr6QIUFgTVcuWLEJLAZfj/tSUDjmPLkkjfIKovv36GFIIIOJ8u1vP9AI25pF
s9uht91yxoxVVJAo55LtlBsuKWIPKmAzwFRlgwOr8k8rx4hRXxpZPMEqGpvaa48S
HrvrItqOevs5TUz51L3OF72d4KSiDqyd+5JLT3qAFY7HipsqJ/LQXQAM6ljM//wy
Jv+WAxBbc5Tx6uRCGrtQJAGYKLQ7Shu8a2r3HAjCQq/84TG59VPD5h1ajcZL8mRt
Gz1kKIjik1nh7msLvtuAsINGXw2lBeubmmvIGl0U8jAm9lQUCFb7lm8QhzL3znT7
oHsikgca6rj99hIE3aDAdjZlysVEgYk/uYoWAG2qerkfzjni5QVfvfa+udqMLR/t
tPWYsZnJ6LC+E80v5lUVUrHLEAHWiWilXCrUze8rBtkwaiwaJXG9SDH6VRj9LdOu
0hNUWrU6ugArb6e2cgRnjChZdPiBZD/DDKJlXQIaWWFdwWydReCvCL8ImwqXfQ5s
Cb/NYkPKiD2/+7Pbo9RMr7JzuiNOO8HMWtFHr+QA7ySmnHfIwn4FmdRjcEVP+Q4l
gAz5HWk0EkX1b5p/5kQOOuMSdQrTMjHsbD7cA9IZRg5vpC7iYcX9nk4PV6dyGLHR
dNMRImxilikvlmXVMJYAKdvEyVzNY8IumNr7F4it4r1YnDxkdzsSV8rcuUWKt/wp
bmTrVNstJfSU0b+Tz4A08NuSVydGa6nsguxdjlXwdBAzLPl6jlAv+gTE1vhmtgB4
txrBQR5bcqoklIw4+m48acwcDINeAS2ZhZXPKu9uircPV8oExCgWy2hLHxymA41R
d8NgCTx7vryTFPfQ0nhuY5sD86+DhBpS5puBdo8xhIIXFmOIsvHaCK6eEC07Vswt
r3cTnu1yIh0MsFIbbs5S+xY84MZz9THCOdw4UbrmahSAK1ZGz9HpP9uDOaHdI+qw
/diMYORPhtGUw7+ljoZy5PEH6p4eHTNOMVPXqik0Zpizkrt9m+EPE6hZYdR1rnz7
2CZeL3YqDmd2LWijCmTW6R8poTHNa1dRnh8YPPKfJ/ctoMNKrvuLSmXmGhaoosBu
fVGXjP501oW6o83CqgEXkwWSfGin3bRSrnSdFjdaaqNh1iMtyWXf5lwKRp3QXEYT
yhXZbo4PIVuw7J8MH4STpFctlPUoCGPl0j8W7o3JM4MPadfbZOWkgd8JNyhALJA8
yHV9f//LNARLTJMZSH5M60LuRUQZxHdQaC3rQBz9T06bLD4BsJCrDUDUCBHjGAtT
Lm22UxoL62brY3mIHis2MvugvW1wzEGBPZve8Llq+U9Yo2gvQTyrMZyuCIkleVIk
qOmWRwi521D4Kf6+NRVvr1yYXV39ZuvFx6Owl2E1wYgM+iTIsMwRLfdJUGPnrAPg
6aBrfRXNF3JwtR9CP9ASjYLp2k3uIuQuHijVZUox1wz4VzLgdbk3O2JZ4KgfYbq7
4nhRXm3bl06WPFP8hYdSd61QwivtjmkOXsGNvUxWLQM66QlooEGoIWCdjkGPnxt3
hVGxTtxune9g1EWLEUpXYNUjIZo+hHvODX2r+TWZraz6BaR+IWgORnWO26v7Nygc
pUSjEZHkR1PKhJyKy6ouEfkFP8Rf9f69UVp/YpP5WA8EeVzSrd6Ih7rvIp9N3kga
rhFPhRzbRdthBPxKLe2ahnLn0Xz01AeN7VcI+cZHAKs8U5Zz5REmvknqtrr+LHxa
BKX5Wz5EnmTnKX4EeyiCsv7EH4e8WSEEk/vnBdZJHIGt82Q1ysWInr4CbNn09qPR
VvOTlpX/3yv9JbLOWqlxr54l4W6io6v/6JB6e0ssn0u237ajj+nA1vOCKTFBq6VO
2erfTtdMvoQ3d/oeJIxeyD8BUMtVLcWq0w0yvIgtAuKyAJ99cbEOcghIBjXVET5z
pBGkSc3XoGRulmmO0uVtslBko+H9nwwcAitwIkR8TExknbFb3PYHa5RltsgAQULA
DI5dEFo3XNvgGAY95/Alu+n6ZkV+k69FE4xMexNAI+/w5kSrwlSJXvr8zeCFqlib
Rj6u6pbehlMy07K/z+ME9k8YICa33bO05qN2D4KeBrJMm2aDAvyxO0sdXeR2yaDJ
YuHmdPNj4dzTsDGBfZ5Ip30A3oLPxnbyqdZ3liH38D8f1kUBwmqdRfeginACWUNN
YhyqsY+XjBFSGIKKYdWVtkZyjbD+5t0963EqXBsCjFJpm7GwtQ7TPjCZv0lN/Vti
tzFhqD/qbnsXNj/SuEflposmj1NydGKCrYCnh0z8jWhSzJcGyMdFZDOqlnsu1rw5
ZeT8jqh5Biv93YFGNA5e9RzLq2JVc0gyC333dSAvn2jTPKEZkXRdygGvZ2gGsqdT
kcWycY1BbC3ZoL3+HIF3QKzLqyRk9vbTgqAddxZvE+5I5ABrGgszNbENiZOlmT63
EriVsXBEV/Xbds0LTa1479Kt35Z0U7TZxnjpuIIisAfsNdh8Obyb6kL7oqHTUcSg
`protect end_protected