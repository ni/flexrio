`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 33072 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
3JbtNiAekMoRUw6FSbjvdAC3OlFvPiEantUwepCKdm7/K87kVtRS/Qbl+d1u3slp
2FcfRSBetTJtJfecwG51nUrLE/TMd396+FDQDxevDF4M0bIqtn7nGORN8psbZlfL
uIRlWWDmHsCJeYb+Emttn6Tbj1CVpdVwO90y/YyV69C5PKUCKlUTF8I5lGnlSE2R
bo0x89qR92I7W9jd0POP+ZYGnEYUcFqmBTpFVo5f6YBtdCqfZl2t+X69fR/sAXvR
kh13duWZNxGfTE1H2YXNedjbheX6GU+hkAT7rV9ZyLxT/mwDDw3yCGWoeSlpajny
9o12lmA0E1Grpsg0zGPbSACQOfKUQ14noRwfGcKyFnXvWkxtmVETiAxAB1NUvQyQ
DlDSULPG3kn4e3+KYiXw/SiF/xqm6BigW/8Cku7GEJVO+GbTGKtM0JnPDxePzk5z
C26v9/eqrlHyvHZjrvz2aLabeJyxwxUt0Xaptvk21wZAmIYNcCTGGvOz6eEvlim3
7Np+dCUft4ZCyxi7NIZm22tvXWpKsFv0MUjuqrYKvDUrzfQROhDCCpoDwu98hKQc
NAVI/Iy/J28x+aIXuw0zWUmMzYTieNinKQEusU0lBnud77+sqWT4dKxtNnoidDbv
66WNcOk1wRqCBfTRl9PLLocH90O2kMmVR2WFi+qhti+RHokdmCOV+8UzmGsoG2Aq
O5BJt1lXBE3v+PyXiJN819hJx69hPDkgSkK0XNEgoSMxkAg/64XOfv3F4gQLQ2fV
BnS+0UsmdDzfNVyM2T3hw6NATMpsXQxZa27WRrW61zaEkhAJFvjf4xPtwXOG8wol
zdxFVNzimfqLKlJKjDz02QjkWJrg6donIhFactMCzqGM/1dm3KaOPONYs175qicJ
4FqyUsF6E8t2pLg9anfzUgiWFxhLZUJwSzcT5XLIkH4/1OjAV5Uja4ZdX/1KdHA6
SoJzJzM7q1hePix/9ouOtTS7X+SwGdyPi2r5h3uItrNdZWRPH8Sv9sspbf4mXpGK
W+XUvvT8kKpW4f1JkjWkgjUDHUx89fZNBYzhOep70YDOdEO9ody2Bizv2XnD/BIQ
YYW4zsXRllVxfuyqQpeVo/1ZIVVt7vkEMoSpmLuPomCtQe+vdMmjKPi8h5wnYNDu
Dr7vb30++cKzCAcLhE6HNGWFB+/LCME1G638ulQc20bvX4qyv9xIhGcdeWLxUZei
Taar0fRg37p6AAXQTYaUCEvF7NDcIejRVHXgj+7buUY6vKvMc8gkCVMnW5rTZisn
78b+3aBNA42qf6k7X/r1KTm3jROFU5Dwks8wTxEsTLAPaOO8H7s/Tt6T2KB0E4AZ
SmId8bq21bSJZRY8k6HSBoZlktNL0eY8PrYQ5bKdslUesiI/yR0InsPPFXG/yF0i
8a58NuqTJCsqE3og2zlfcpQxA1uqKTT9TQmRBAssKBeflkxi0XVLLMN4rC04hoGA
S4j3DuSX4ppkXGBcIe3CRdpM1NulAObkhh7h8eRDoL3MPGsVHFHbIz3wGDs88PKX
8tOkeZWUyCz7w0pc5gUZDOz1PDUsWm+PuXQmquYIUiW+Y+AGd89Iwk1hKgX3VMIm
5PFdTUw9y2wrn1j2QehudZf8hdwfcubOlwSuSzJ3+Mk4QINFxuYa4V/n3xtzx8MK
fRw7Z4oKEC+dvvJFEaSsjXW9pWShA3J73tx/m2iDm1gOrVHoKKZnEXIC56IlVL8R
t5Vismrd8HoQpm5r24saVtRUJ/0J34NAU9t1+imQFsjbGpZY9SA+HlUnLv9TAAo5
KZYmyHPq3wx0q2oMF/Pp45PT0+mqG4BoY0SMmIjAzHG4S332ARk4k84izwT7Lh3S
x5k0rRzbCxadR2UAwt7StkKdWMgJHCvC9lvljuFUzyQ74VVPGlQcHznYVpuEvG8L
YwbfeWu9wPuQlhX4oD16XqA6XtyXc63Cyf8059rIGnwqrSRZ7n1knJ2ZupHTdmCx
sWOvUeYfgVTKB8Qc93UKYmdwN2FL14ZzbXoLv3BkZUcXr9DQl6kVzOpzn3qdaZMQ
gn3Quq5r0wbdZ2xMl0U9RbjMcz5+g7lepk5mmPd1RHBckE8WSHvbQ6zkdsfsgoI9
DsCIe7Zf9SywOQEfVamanalOYJvsX1crBe5/cqix5XMyaWz3VmeihOX6wgfoZTcF
O2bVrQRoQswbxAciio7fMsG1wMwpx+pzrWBtzgtaRuHafR7tYsBalm/s5G4cayrq
5q/J7Q20t8542f0cwCE/jxqLp+7Px2RpJwE84VgLMXLY9UHOMo7y2cKQrjtfwC2R
v48dENKdvqN9R87IpTUWl1mvAQAW7N/Pawg37Uv2lFb9NBhFGCP9SSy84i1hiIau
Tksgxpkn3Kq61smcxwOwxokIrgDzaUSePSfIx83DDotWus70sd+5YugblAtbWgyF
RHp40JbV8rzDAc1eVAREUrXMM7zMJrPPqrBBurDAun9as0VEk7fXOwYhZVSkY+Xs
HOUqbYDarVfmzbcMp+/M3xULUJjQv7UpwH07UP0Rq/NMOg/tLW4oM12H4mBE//51
vEDluirU/l5jkjenoC/k/ZeR0nBHPFaDhx6MD5aPZrvI7qDBCEyzJbvCRNp51rtE
5A8NFThdOaTASRRv+PNGzG3Ffm84SxC6KEM+ZARbu+k+JLcS+KYZ12nXk1xxPtb0
bUu3jzN9mizJMpkHZCqV4Fv4ZYIG/39xZyv9ZQUL+PFi36O8b/f9ncw5As6C7ldz
sTEUZB5TqARc4hFglo8fv5MDvTREH5cLcc49krPZdsYa0B90cGRVHEj6uWNGQIez
w4ZD+y0dceOZeYutF03TRiEmzxGLy5QKn6h6zm4/G++U96MiEMjDhoR2wYlniNsq
7mts/7nAkqIxGxTZLM/1/TQUOYjFga3rqqBnVAPFbKdaX4ztI8LqE8iZUQhk0low
vpoOQ4SmMjq+p6ia6T+3/CekGD7rc+1w3YKLtfLCyTQlLduoLajjlJ0K11hcvQml
S0lPzzELNe4QgyCFoDOwRmBY5TQOg6P73ukV1tJD/681HuQngeKQpgKoc07twiu5
32DatSBvybKBcLh8pagpmcv7qKPuF2immQKKfyUXzONMqm8mzemcJLkf+eyXhXLG
2UDr+wHMB00xk6rEi/bH6DtXCVmNW+74TEZUZKUfUeot5JnaadMx+8rd5BF5yTkx
fJcsd+r4WzGv4rgqyVlZBQ0WIog2mIYM3uJre11xPxgtu1PvclSWTPTb+x6kozmq
Sy4Ej/Tbs+7Y5F9gCf1cAZ6XXPI6JyJK8N8KMlEm7Gp/MOf5Q5ueDmIzruC4i7Hg
vt9JdOOQ3fgPQSNY1O5iS0iG/StNyOB+2ekNzjxcxsriTxD+mXc6MezPhzPzr+JQ
bwjWTOiSbyIT8+acMCTL0rMhy6dO02ph56VuWdNn9IGq02EsubJDAIAr4SoyVYEY
q3VBdt6BzPYckpWbO8sxghzXPrDhOMRs3HjVYxW5EERJ7OwVuN4f3+t/XvOY3W7K
0+dXH8IA0re0raJ+3Du35shnBCunZuZmGPNAqOwiALDg6eKaFvdhegjDZ2MkDWxB
5U5Z8/mK99F7UplWkRFe9ncIyDJBgB5IlT8wDGYfedLfGBXY8/n8FH77833Il+Jw
pq5VZWBTylregLyy8n9K0M0JHZDBUlJcvCmrm08ehaTpmbxXeQKg6/utNPKus+se
KrE4kdbSZJ8izjnic77hO6nvDYIvDWYc5QcObWKtJzAX0wn4vJibXMwCIoFyH1Pf
tNRux0oD8R36LheYhLEUIV+NVl/1omTJe0JU2dpTaHTUMmOPNWc+kMz/tuAFrNwC
Icshs/epL9yragZy94M4ADZoGqWN9y6E0GBrTHsoho3Mubh1vMoXGdr3SKpJqlpN
ntM66iVYFFnPwxBLyuevrE+VZFrzXIVI1v0Lp+03XJm2f1ZQn6CenIGR+VauhEMc
PaaclRgXoTiUfCW73+y1GdJB8heQiPNnG2GVLIjw9BdcZ9lF26k1YPcTqiMhmBwx
IkoRzG392DEfhDSQiGjUAGu6l9aWlLW8Gggx/2Ud4BLQnKkzw1rpR1CorfB++Mc2
ZGH9JxYXAWzVccLx2w/eRtXIXN0JPPb5Mfh0YGv/BpDqFZADBCvG3x7wUsqApxmI
4BGvy7ZzEuuSUwzVSXWnz3rmLRRVwMJcecT8engAEUJEyiH2Sk9CMjv0rqB5nWlA
/aF8bF9JOk9Em8wI8c8ls/HQ66z66JNqwWa+doVgPHC1FbBZXwPVLn7nYbLEPi3E
aD++fzWu28n8BKeqNJQe3mI/te8rWExChPDVhizcY3oT38N7gcP7aU0rCZ0ueuE7
EkwJaEUcaMa2heUY1C9Y6TwTBsiap5MewanBYxiBxh9LkMDmE9kOZ2TIStD1T9H8
TmmcHBEL0YhKHgo2rdnyXJR+WwAW0lFVnvZjO1zN2EN6+lztbTHz336FIOINxxry
v8lBiQLOAYXkXRJP1Kv44x4VPsPwt9Y4W2ph97gP2jETSMF8c+QFdaJFMhybO1y0
pe9XboISwGS6s1nKLv7nRyIcTJO5ETiwiSiEAbF8KwCZtII1/l62db114JPUFUlZ
T26Ry4TpgJLHCLbsb22jcUNZfKsPtPMUbAhOAz9IgzkH7abRPjowbo9MiEprm+e8
/aNjnnfyrNFvvOVSo3wWHOsW8gq5tY21ACT1SHPAUWMdmTsowBnIfSUr7fCDbpb5
QE+OEdSAqr6LYMibhRyG9P6bYdkjKnaPRK8/bWrD8UCdgm7cZR5hteItDJSi0tRN
GNFGxdtgoEqE+P1PV7P3c6LZkX+cKJZkAVckNdHA/TEtGHzY1P/e5oEZ2YA+qMOi
AW4qJwTKfOV5jNecm+29fEUIkNqFwfG1cuw4N421NNciiPDIR2K+uTn6BF6SBsYU
SXswd0MxDHWd+7B/7Bvp1maes9pBdrQu24RehGvnra5m4wFBadh/T3mgY1dfmCj0
+gDw0B3IiYIu15vzo/nj32ywIaDGFvmUSlfJy6mZ+oNhIAco5hjHVjCQM+zjPk+o
TQGQyGko0DZpTZhuA6sXVfVg7iMBlaBLLSv7rDBn9dE2QLIv67YAcj+nGFF0groH
bt5makaElZmVLwix6lxHzs0+LvyytR9SFMGZ/IJfUGeUHUNfttjxEc7OqIIwKqAY
g8sW6QoWOIxUQex1cbVyPALgFRgtw8SSQqlz9VXn9k5p7QUIciuSRQZr2tOkUpO5
+OTGBWU04xaaZaOKI7DGP8S9mtptR9D2HSgwLr/NsQU+8LX0M0bemdf2R1WAnmZz
sUr9KC0toYbVGgrTb0r8Xbr8Wlsjyeyw3u6wWMOFvQXoaX26ctNbbvSzUpbaVrnU
7e+Sj8bB8FAUvBQeGcve41fvHNa/Vt2iCGmM8PDyFogQV58vgtp45LpwHbSwJvCa
2QY8vKQXjgNbuumB99thf5LUVSl2QQeoPal6Npy9/lCLwAID7LucN8mUHYEjS1r9
dXv44HID7P4JvhREMZFvtKjNKJbNWcRlIeNZgQ1G8zIBcDykW3es80xT5BUx7l3c
lOgiiufMOox1/3la/XNKE4b/HQIcgYXseeKVYnTZtHbSEr5xT7RVEzevd7uWIBK8
rMKcjQbcWa/kGiRW2gdpm/OJzDQneHlE2v9JOKqib54sx9DYcpA3wb58FbWArGxp
ZgrkO02IfwaMyaQpLjgCmFy17GFIeTgeYShN6dKLJ0yG7zm7ZC0WJnuGnXFrURRQ
0hXNUEGPW9l2Ha3qMDvzDcVURwgA4RvxuyJ26ENpyNj+BzFe1iu/cw3GORdAUqCQ
n7e0mo9+zJ6ek0TJW961e7WsLB3iF6a+NxFrM5LFEj9TnVl39qYXM49AzRF7SK7y
EMpZNYomGj2dYUOmkpKezw5vkSYd2DWqXeVYspc+bu3sdbhPUPWAWwVK+7ZNm8Gl
DRNHyrRkuDEIqWPKJI7Q6Kx+CGlBBpiQF1oYoYKkwd4/7h58UgEZxCHcZS/xXYg0
wC1O1/KMH41SSzutZ7pEGtOks4+IDgyL7xLgYoq5HEbUWG2bO5gBoxWN4sJPvvC8
JGQTDb8E4reUr06YUvhCrFbV6boiwVglUdGwXIeAFFUgzfVlx8enIn+H+uby9wdp
S5HRetBKbRa9syZk+0PyKQTSVbZX8pXR45ZIoekDlrGYMObpJbDZkyVjwQ3yqAAB
fT4xl+p0yTkt1exzonPHbOiWRQKD4Vi/nGMeSC9GRI+0ipVlHa3yl7pbqeZXJ6yw
pHL6PqilxNq8iCShKt/cG4cKVsVgri73HZj3zDX0jVrSW5JogAu8lz9eaxH8v+lP
ijHhnpCqnhLS+UBsFc3RAryKfYopjcJ2mz07TTZPc5WPy/Cx+H65ohIlGIBQcYRm
5ZPq0i9KqHfZTvIrDhg757BjKYyKR0tCwEUCRBwUFKWW3KAAFXC2Cl9DGHZn1BsX
U6dLpWiVlydRbupx4t1QsKdYwY0Tf8uH4rQR5EjrpyUWeX9pExpCyli3YDQOrLXN
FGXzMVvuYe7vPlUfqP/1jnzzdw0HlpGy439U7b7uIgtUDwXXoVnkVbOITuUoIBja
6jm/N9zEE5/PL+1I8hNcwQYGWBPMwSRF9GYn0X+zXPCG+WQMfiT5w0Nad8nGwDaE
7GaUIR6JaVMDTS2tG41Xg5iavhUQF71thk2J1tbZroje4Fwd3TT3M82kpPGPE5RG
xHQ5QDaxrrzoaMTgeSKpeSCo9sjuoQs9YkGRuiXCO4ALgYt0MiFOCROdLVEeBEIr
z00H/6/8zByZEy1aeUPRj10OxOKdWIZnSwko3qNj2grggejF7EpFTZdEL1R6bDHd
noZsjkiu7TPSO97zNMZfv6+Xm0GoLm8cSsaGbX2gldDIX6bT/3F8ZZ8w3X/mBDEs
u1ODb091YkPw0IGAWJj9FZl2vTBqpvw/W3mpMWlh9j2Qp3OawlgUJZkvGBBingDh
DpjKQCHNnb/ymFg/YyKe97u84KwKz1e4sBH6CSzP9QpuB0x6PRtdnn4FhEbCjFSo
a05ISayrdo9E/fMwvDhKtD7/VE5JY9GuH+y7gfeTifF69s+0ObXjhOCCHyRFnvvb
1uCK7yyPdyYeDOEaqhMgauf9nt3ehDysNnjXyieWkXgMXwuPMTg445YbYVxB3cUc
CAsD9ZFNUnUS2EusefvxBny949ZUC0JycVBvm/p4xnZNSttDHJGOjvEFvbfjyhtp
esQhdvKyZXfRPvbJEN5LeFByRYskHQfl59ZpQgs0gd366UkMorzRZCMofGYADrV9
xM8fJ0wqxalzmKpLoebEh4+lIU1g6d0m1iaLbNLkDBoSEnU4QeHI5J4zeiiEpUr2
Fgj0mcsJCxe1E5mj0hmXbbE4CB1VwhaA8fSuMvf74Na5AZHSt4wZV+MNebaxPNSL
gL8geNTM8ytcB8s0YGyfAraLgiDj4VYleBb+JskxnYOIJOwttzNTIYKXthlbWHLT
gNE+Ok60N3ZWH2YTejyKtt7UbgU09LndHJBr1yUpUl6FFkilhKPhXzx+wykyscwc
/D1hrMhbAkmB9SKUS7AljFJpHbfmiPQ5/KPZOiwexpL5ccF1CkJvG5iI0erMCbzL
fv1Xc7vdkFeo1r1uKY+e2sKuxprWZqbad30oFM6N0wQBWKeNDLIOySyzNvFNCgD4
V9diUUyL3heR8M1jV54Xr1fz1aUlwtl/dUN/bWSjOUEj+Y/xMBPAKUuvBpb3YB/k
PqePiJaeIFaK9xn+DaduLlR9VCNyZ+nS8gjKTClWMnkGYOH9QSyXFZlEg8aV0JMG
X8/leEmQMi9K5P51N52HTkmI1q3IqVKJpUb0dBcCT7MUkH7Z06AVl+4soVyWs2oy
/4x3U8LDJ/LLM2srEVV0fuVjisu2F6h/lSicnpMsgQnJ/EGLCnLmaT8TZwZxHWIX
QprilYJ6VgW7S6TZ2cCz+5A1Pa8bdfX8fhJkoo5dFDtjukTZaVPi1sIwDMZL77Gb
HahvgoA7WbNFN57ww1p7haE8OLGV/xDUQf3kPDf8f3XpWBRgCxUUhGYnHLPVAJzj
gLv952q/3/3XjH2Gb6jqFPm/hIf3feco2B8rDn/IhjPnX3+C1QoTQgzwbQniMraz
8IBQHUmRlEBZnLqxf/3K5Mjqv2/ESLQkvq4hO/guVPNACJddpeY+J/tgXa6M4P8e
aDjitERgr2HCGezEywvlYvhYJNyNKYV/7eJ5uMbz+UuSBmQp9OpZFllvbZkTuDY5
BC54iCuAm/+0B089hdQGxOuRKen+Y3sx8OqPDzUOiJcp40uNZ+pFanyyWfDpV4ds
1QGTNhLC8k+24dlZsbHH+4lT2kO/c4EVRVD2/6HCo44bsnFBDWUjytnyp7n0+dei
JylbFBQ+ScVyJkk03DzRyPUDyUbdety0/lOFEBOpQF6arOdzaIK8TJsbtpgBUujh
4DkBTvuSYd3urymSB2iApLCgrr7sLVbgdb0IxoQooMoR1roMdVvCmhGMUIJqC1Fj
kE7e+WiuDA6VRtEtGqXGoV+A4EP6A6RNUpQqXecXSeHwn+xvLk3XH3ZhPgvSadMG
geGsgAe09KxdvS/dIu4rIxp4G3se9iONCHDb0pktKMcGMhFbLfb0Rp/HBWD8Wy8I
4azea/WyTcfFi/+a8ULiVU3C4+dglafn2BFhwk5MbedvIRgH4ZK3mR1cbNNENPe8
OuOKfZzYwC5qtcboGIBOCni9IFX6tYb3tPfx22pRhFbetTMdy/Jj9quMsT4jcxCr
1A/Gfr7AMBcB6uqNnOwA1xqoyCN2DuIYjL0Du7oEwOhYs8pjhOhAcqhSSLSj5ZdJ
hI5bemOpx7Kiabur6UIpB91oXcZ7ouUdiGLqU+7RkSyBOAW/LrtTCccDOQdJAW+y
t0KLN8EuG5jfCkrxVDwpNRwWhv1ZFubK2bBjTvEzqgT9kFauwPZ0msamx2xi2bku
BeDadfiyhGeB2GQKWEECntkt31hRNfyRMlhbOOa6HzBeto3WFW+90mmwkWeHXv6Y
Dw0iafFNZX9B/W1DcSHCeS7bGeNxUG/+UwMCnh2dlWsnQG4uMrJ+ZIcFNWb6YLnC
gwsqxAWmHZPoPQ/9N+sk0hoAxyYbm/rRQpCf4fB53c5+DQVFCphp4NZ4zFve4mVN
zVtGe1cTkBPzywq2fevpL+8IWKJBrM8Z1xJk6pC53t7+ql4+PBJYcrCb3cYvs6cO
8+5m0SkzruxM0fTq2I3n6GmQ81apCr8MXTFK35FUMn01eXCTV8Mj+UKS8fFNVC1k
jtjOLKIFwIGWwMZDqOiwnM10otr2Y1v6i+6wQl2ttSyhkmFVQg9xm5+Few6dbbyj
u1d3q1q/y6tGKoHzxbkQMmVepzk5rrO4Bf+sVbrPF7ArIrCwZPLvfJP0i0TCmtMw
pNEnPeD+NwLn/znXFoflLuPKUDe85bA303XDcGA8Fj/lP1ZpesG6HFkp/DArEivo
ywU9dDaQzAT2ocJzYkLZhWLuLtc+4dcYMXoy+r6e/U8p5miRXRZuzMHbLuk40yl+
TMrnwfhrZKubvAD+/BdPQZofKlkeWWbs8mRejqg974HDGc5FHfc1P/nILRwG3l4T
HFRgS6DokE7ZuUIKTeqAZznv0l7nt57fkHYx24nKIR/y0IB9GsOdWnh3hsiLPoLv
85VRgRKppGMxO8LkkfXdPVu8RMQLzx4uooka7cvKTunHp8TDH7DIH4UeEEZ1bzDI
LGPj5IVO5rzOR4Ck+UVoDL7+5vJHTj9JvCPa7VaezeVMzDGrEsIX/0Dou2VeK5Yh
GmQoN53bJqDiecHN0p4bvRDp9dxiRw0kyePxKvy3w/VHwvcr52i+aA9cDuw2bZnZ
qazRpN4GoTB7m04eHIvim6a1z1z+LfrEfkEbG9oB8bGzBNzb+NS5LPHXdwQecKPM
cP024/1x9D4lsLUAAk5f5CyMzXKQuOdkEIZZjBKjpFRDOfTaELBboA7r9O36M9s7
hEPCq4u/Af9YYJnks7VaFsTGjyrUoEHpmZyl3l7ffLnbKgnx5Z2ELshxjhIGp2zT
MVh0dGCksgPVgAXA4z/RyLWia1Ds9MTd+KCjviTr6m26Sq+5gU0F3ZjIky4bdhya
uiEyyJ3zAWJdxOCipN7z62pYpaiPZic/ixa45H0aqEsVwWIr7uynvTu5PUlPDw9+
afLnJS7WmzlcAT6eWt0JUC9oOtAePt1rnC/ar0Yw2AVHZUDjzCN/7b6mXm714Qy1
AshOK9FXrFMt2ZmtedvDwP+vErj5TkkFk108FkGm6sjW6lFVhkkwpKOlAf7H6Pa7
jJdh9Cd3zQ5aggjRJDI++VKJTv+6XA5+YF5I2p/EUqUSIpTSKHzrfayLO1kQJQfL
IVdtGiJfim5ElJg/RT5tM5EY7yuJ0rPyO4yaigl8O/ba7Adb0LaAwDyepl8VZJEI
sCb5cIcTwkyljaroEP4P2GxVfsmnG79gXMeXQeOWYZnmMqKz5jzz5TT7UziPI0WO
USW1ub4cCDQr38GbjphM+UHjTrZhsXMsxFfX3oVgP/RkINwsw0O9pUPQzvhHUcB7
gnfP32jqxfz4ypTtUpY70UoWFIvN8XmWIfk99t07c2Pgm8CfOhy39GHZSx3qKhzf
OlwR4Ac3zyB7t3Bga0zPavLiimYjiREWgRLSd4k2pWXKtVifpSsJCCC6GPP0GfgW
o2qmGJUDVT+5pHhZmjB/bKREQox8myn2RY4jehLqIsaRQIaiG89qc7gZTdpButHc
r4/+7gCh8U4YCoFrDFIZAVxr6NHjzPAdcjQexwSUc/8A5saw/hH3WxhizkVHwg1s
7OLv52QSekpnyXFtrFZ8kGUM8nZlejrYgKhdZVrkr8TpnWdmRhQxrnD5MyBvd7R1
yPdG9z2xpCZGRxzBwdjbDYGA/xrAImLC8gs64RVjLxomyfAcsStvn3w3g2fPjMqp
rn9YumA0b9KGW+M0K706jsdp/hd2FDWzTenl4zDcl/ti0N2L1HBfIvsLOpQWusDR
xKVUQAM1jhCxO5kgYEkqLVcX1ALOAE3+ufJJhGM8mY8WXmayWtlTNtwNnvCWtH6i
Tm34uUIogPW8ZAm7C5dWRqkibWckj31S9TVpEyJCIE200A0GdxjRbfA/12iJFcqv
NGbz37eLd5AsVTG3IAfwUbYh3IFC0fSnnH9SBBiUTB2uIxItEWh8UcgiqLT9WeH+
lBZieJGNH++04UC+2UEXNn+tG0dTYc8ZBwTJBKS104n9ZLSFtcbKdJcJMVwlql7j
3wSFXhFqoLF8Izk3T56/zy3yHgQ1ZoPP4+mavFYCqhKGgwRY9x8ujAX7ui57jaqC
KSVqOS62eybT0NhSXwLO8m+OuI+IgUDOGMXBsd35ZuFdCQLZqTpmTiTTNefEDtcz
D669JQegwrJOa+fgcSlfymVsM3Ws3k+xoGPjgPvIlUfwgCTp0hVB/7F7S9feuEzw
PQDgC3b+aNDawN4Igdq8qS3RNRtfx9QXriecKoh29leCoN5LbxzaL/PlwuWhovec
lSwNgTTj/kinrGbz7PDhVuGBiOEogsCGIl6aeDXs+Ak5SD8KWvGKxnIB5x8w3jnA
q5DXKR/CXiI/3felgpTHpZARyPTykUVptegPtkeNEfu0rgBOeVVZaa/LNFD7pUME
41ptizIXVGRJ9EbNkGVicqjg7kWq0C8FiSMoZXNz09N6I7WizYOXekFjRepzCVWh
Hh0WZ/0yJN+MWX5N41BFgorguTR++4gsXNB1W71xrQb00SuJ2LRAg03jzJOTOAs/
l9QaM+L8RiRu9ScOq3CgyY6f3R3TduNWXKASSjCN+eCqhY2rsaHXA8jkGbP1Z9uU
9ZO3Y35dxg8YAD5rXY6LEHAw3FHA1S9lZK6nd3vlJqmGA4+9sCpeWS3UHGYdn27c
B6hHWB2x2NMLgfC6pg7rHgZncnzRyQnDjSopLnzPDJAG2/AbBIlfrLCpeM8wLlgx
aDe2rAa1nDzrg2qdLqHua35iERvX7fZfNApmwNWY0zwPSKIctntaL2kJrK6nMS4o
NvaIi3mYekhqMzNGJx7rVD7QtHbPneuKkzmTNh9/pdwA/0bjmLtBxYauALMYEDCQ
9zgKn3ZWHlIwDkz5eLpxkeY8Cfoz9dbLcIqS6hCdlsUe35hOswPDre/w4w+2bn/C
Klyp6NgMe6K5h97BFi7grIjrsdXP4n+CMIIOximBdztcy28N/tZT6p1fjc+6zIYM
Yyobl+4iRNnijPVF+zzYbns82T/Xm3lDjQuN2jKlkQHYE1gi/fvnQ4VBJg4Hq5Ew
TJltE1MVe4LI9k/fqsRHMtSatYzNt7TQOXRpeO07tsB10OQg+NY6sTYX4EBcU1i4
/avIXcXmuI+Bl2yXcSjaaHmnCl5Yi5YVjNN2RI0yc69mB/Ufz6PXUuVC5BSc0JLv
vZEc/mv9GhVjh1kvkee40NqOgyylLF3dTrcGW/TJ6I/MgqxxgELQYU9ZjvJ1t1ii
if/zhIGXvxnDSnqdkg3b6diHKV5VQaAmGk0wuj5ENhbcAub/FQgSHNOBiDDHNTwF
Ox3ru3NKD6dGszFUPlvc20DbNX7o9Ce7FpJy/FxGq+hQxQ6GTyqBrPqQCN8asVpj
iRp/V483bngtDPafcyO6z3zCVu152uGVpNXMwoOuvpDcBKYEO/GTdaOo6Q6FgBI9
8bxmJ/Gtr5xhPX+dGe0tZhdDxA20rxEisrZ1eiYNIFLeyN4njNJpEpW7Q/MwIHjI
sL9iidXysBj8noB99ohdRtdp0LUu4gZ9ZoKMKREWnlSw04necD//8N71ByTm2tCL
jKVkqMGvbFB1OzYPzvqMYvzOvoEFJ+dKDqZa8eT4fsmxKRrfrwNOn39nnppdPZAU
28yUG9HDCydTpsCclyYgoC380wH05LU6WIKSad11YfAJYymtGaJPUjbsuA9/0/Nr
UybUs4vlBqM16B5sQfk6lUmjIUiThfZdgQd12118IhR3XhghI4dBk6oP7ekPVAWf
+RcIjrPfKLASH/Y+SPkCWLPfMKipJFcnVkThL89X6yFRW4ho+5l+VyO+q8m7+2wS
EXsHeaxiaH3DYI54DpVvvAuZI6TIiAx7MKxn3/ET9ThwH6wK/txJYLTzEYvaXH6t
OsrTDIyQHG0nLPCy1cVzM8udyUQuBQx5CG80akVKgI6WIi+/6Dl8v9ZJinFsNiqh
jAX5Qkqy6K/GwTOxLs+edLDbAIcjIOVe2ujr89IynFgb/9jvPEX7z8EyHMyz8Sw/
IKlA6U3Pw1bKa5xkJuwfE5qWMZqUAhEyRaqFifdB+0imgQ8BMyc+Y+H6O8OuaJ4w
8oP4lVdf/DWbBKer2tfyuNbKyaYCoW/K7FTeFrhAvoTLnMjy02g52vTjHoB+EA/B
x3Zhq6WJZ3Q8wfZz8c2Z8dmnEVpOH9dxLP5VPrzj5y9QB9AhdcBLnF9Od0kn0W7M
jpBowS8ABAzu8utHop9vVRUkewuV36T0XC+7KAfAA5u01ed+gCANu/Q/ZWVOWNfA
XCh7OpdRFmIhePbQevKtRfyH+y1Vwl0kw62Q/sp5SZXhkm+ZUvv9xXGsbHyvRRAn
7ndxaM9bkU6ojf3uuGYgXxzAiM/VxA+KkEgr7EUpxnVaJizJ0e0KNN/dT2npCpKN
NnCvQp/+2mGm8SCg2iC5576JDeAF5rIw6DG87DmHX+cKwWGkdtbiA0VVfZyKMHsM
PTw4dDtRU0winZfJUAiUdZJtSAlGUCFfaJOihCwlzm26gXd3qdsJKr9RVq9zC2XY
QDgeysB65AGeCU5T+8lwysCXpnxOvc748YFXQdZ3WjgMivfaZylH8Pr+s0R+43ua
UNPaFZ//i4Amu/BxHa60PQa4VCkm8IOx0m8u24w6OVnbu2TyKH7gatsyPVFcTESN
G9N4yOgD8Tz0jpBE8+u0aTBgrfKv7BIAKQEN9h7jP8y2XmAMHOc9/aeFJ3b/pMEq
SoW9qIhsiXx80fbKqPEeRfkc540GU9GGFmH0G1CSSLk7P7Uf9601E+xFgAdhJUrP
xpEuNtCyzvuacuzOhil6e2k2qaZUIsn5HBRjv0cY5VJhzJ9vS8uczeHrSXYdlOFV
Q7w2ukcZRG+2z1L1imH6/YwYQdFp7cFhJod+VxdxxFt5UimD8Q+TdomVdsnBHuGN
RgGe62rkStEToeOxfglHHr7u80ABtZ64Ll+q/UQivoIAqGtjx5o/RJD3yTQi5gvk
pLZz6YTAYT72/a/20yLDz1U59QPzgE58tfAw9Pi/hsPehyvzdyDBtcOEo7qQNngg
V6tTfWWh70xeTOpwMd3Etoh0Fv5T6JehMjHtGxjfEZ4j3qz4jkAOV5FksfoJCDSj
Z9XpYMB1RKuULSx7XKEq3nwFA9fJN0t4Q0GCnHv3UPGtEJlUV7hSneXRGtT/a7F0
6Dx8MEdQvO9+MZwh/zla1sM9FwMd0eYOK6mbxMLDKldGjQXhMoYN4Tn6FEMf/7e+
bITq63NBn6ZJ2eebu4P5mUld+vHJZCXeYtwpqz8AYt1Vi8O4MxC1blUsdWr3RQfM
VXhts6TmYARvzCe+NkIfQp/klzytQ7C0LKf1fZvVTuN5fMKFATN88VNMRfTPE/LO
fJECip5DGvO/M1ncK3oS/gK/b9u2tVLXiiegQlQ9vcrxbd8hF3kQoPiSR0G4MA49
Z1bhpvod99Lg0Rzt9walckr6+vpsOrrSYgWlEqc8tp1o7gEZwTJzfjatiZtAHOl1
RjTlR5+fut9TGDbfZkkTN+/HmDG39MD8nBGi0rToHwV0VNe2mxw94G7zOpiSefca
uFuyWvXt0vBCP4rzDIIt17sXICn0mSeDrsS7tAk9RPe6BFLafypvXz9lHgMv0P5E
62bQGxKp42T/ez+Vv/hupeVGKK+AvEOXd3yvmsueDXsJWJbAq08le3IowehK2v7B
EcPzzQESbSt5DVTs9Wo2esJNR9vk9siy7u05TI/Wc+Mz4CbjifAWi6XHTDH1Kljd
TDIyJVXxVsm4nfVdpcMeowfsZGcoNP3d/Q0qN4ewZB6fnp/hM/EfB17greusuZTG
jj07pSB6LhOcy7zLJ/yq6WgRGqULUxcr4Tm1LyE6P/l2S8zyHnDgBn4tBz0BaTE2
+O2LMtd/SmwJfyYibMvsJowP516/TYxwnsRHR1UKBP+zikwxlZHNQgHr+ifsRnHs
KYWbQEIyYWCX/OkazaaGNoPOh1xEG5QRpWg7cabXDW8NldRDmLhi+xYmAxVfaY8i
DCBJsMxGXHEIWrIg4Vdgw+TmO5/VT2JUk87LHpHO4WV26NZ/CdFMWcRD1GrqkOpZ
xaFDXsD66Fiwf2rp6MqyUDB8KDm5fXjPrtAs+q7CO6I+RVc7Ws+nuTTGTdTQkfwt
bMpjDw56lymQkW5BnQkIZHNztsqKDC0gHOINygA6XGrUc+83mzybSCUjcR3h5RCl
de1NQ1v+dNgFhIpQtmkWqDpy6K0y/PQCrEPtltklkjtuJDBHon0iNN8XEII55Z2j
dLGJXEpNSKYtZt5w2EKfAQZqdLwUwkdGetrDZ9V26TczN2nB3prtgJqvLUYwUGak
z02qIS/gqBZN2DI4OdGFYIBTOmeBbNrb8g1eT/kVA7524TD6LwTA1piENv0kMaQm
6I/Cbnk/hBI+UqJO2u1B9as1dMm1QGpzkJA4VctcduPy4LwIhUbSvXPWBqge2ljO
jq+VDmqTCGYsQYDoE/AjiJQGgSJBXJ43YsJJxyqeWC2vJFj033xbeN4j0fqRZCm0
mIqVmksZ5rlCVwIYrhuWKTKACRKqqXtAyBNuafGR8QSLFRk2dX9o2IWVFNk8XlkJ
sVda+0qwoDe799rGGJeMLatgG9x1xmbvpDKL+BX/a+Pj4BJg43veGqq3beU5Znud
w3jkV+UktpXJmppaOb9FSdr4ub4zGbGadpGwjbXK7sTr9fDDwQmhhn5hbvnldTlp
BI0jkjNvOToDv3vL0AB+NTPLahIFiZuvq4XrcrCBT7MrFy9O/fAoV9r9VEZYq43S
28axLdr9Qc0Cx8g9tH5DjLpV+qT68Pd2vUxktnGH43AyVexbhW0CAP4v0pUp6ryF
tMnJ7WScmDqjFKTRkJrp2YEvUzyQxQh7UpXBfV9vj6iOCil7bnzeXnecAPTgLJzc
ylpqlbwpDKwJu1aNo9nE1fB433RLnaRopoVfyHHUubKdr6sKS+uAGZ37LbwHWfRJ
cwwC6wwPBz9bsGSNJ0KNjg3qwX5tZLsdtxRZH1T3kfW2AEpVDQe4gj4OwgUh5LJb
mf1ROkdP64OdViW3itwMoPkgrsyzaGrgVUo54P7RtF72N5+5HAeeeOnDFn629Eqj
ZyWggQ6L/4/N9i5aCOxzLL16j2trSnrjI7aBe2m2HRKTsUWRx+MxP30Y3oX5CdKj
MQVzGykxczcZC6p36QNV9/BBm0JhcUTYZZzjJUfGBeMAOYOmmXTbbGDwF2OX1rkw
1QpTR8YCr1vvpGTv71Q7Um0Mg88WCNlvmCe5LD8NWBHi+vLMQ1YyEeLPueai9FNx
hDzY2h0JW3gCAkkg/JD2n6NWyWb7MCzSIAQ5n3D0oRiENS9HeGH3swyQeJSyYM5i
p+6Zqdi0pAw3lzyTV9bi6F27qHEH+BX2NPvzqmqkzexdaNmPEmgBSI8AA5B2LKUO
zt6oz0vqVS4hJjXNoH9BnHaxTdqqoaPPgJnkUd/lyNdnAqWeCz5qUeVpvq28DlHa
J7sBKop5Y+h3be7a44bCd71x5R6X3OQCgY0Y2JOrWMjuGrTf0WSa0QlBpImXwbOR
JagXkG0tCFxIqKvc+XoO0oqB/3nSMSGAYfdH62C3c2TRGdmmgseTW8FUiTxs14JM
HnVap6p21dUIqdk8aTGgT8SfV5CYwXyczRq8xkQQq4sIwxIkNvQ8MOvw8Ikj4whM
3Be0vW3h/oEPlTNSIcOfuMLZwbibLPzgDx1BPDJAUAtKxMw0K3ULMAFxFPsST7Gr
RttiKcD7pjPXwKZcuOWkAbV26Nlb0ooWSam45W3FE6wf6ywTmAMo/IkDFg/tlj+R
OwXFTQZ3xivlVW0ITEoww5LtJb5gyM2cyF+tuPwmJGtVOeK29fvt7mFCuKoufpAI
xry+log+4lxuEb9wEZbNGpGEStbmEM3eZnqI/jpY//eYHWRoS4GxkNtglHkmWkGK
dt1/l3PoxlkGI1JOXRY2lzV25Ptp3OlwQGjj4E9z6xeyUucVS5wsSV0r3aQybb3v
8WV44EuoiMr/221SkwD24KQcdZ7mF/ZA6CnBWAv3+SBA1bR4bPqj2e2awssg+nbV
k5F0JNAVSQ5Bk44Mgp1VIJVpraut3CUNGp4CRiLUt9Uh3jzBa050gDz4MZsoR7h/
yQvZOLssniilXnNj9pTRJjp1Xqxkt3o2XkF9gJbn1iuKcqpGFx+9v3SpNaI1MbRd
04GDfnEcuonbZcw+MlyKrerXWqIfcnYcGy2DAHEAHj5HQnCp1TfpSoRpef//3i9X
KSdFjNginAgMs1i7Ex7e1a2t/N0o3MQnjK5VdBsGGAf0xCkv9LMHDo3RMDDmJ0cA
nAAOsAFDbyTmxb7PQTOr3InSMe2G0LEPYub+Uv7HlMrjZn+cLqA+4sRAvVgZziO4
j7L/i1pReXh99Fxm3vGnwIvaMgk+5OY93INrO3NPcU325GcZSqo2SJHDOUhBNCjv
ZVlEdy8rXdO+Sj4jDg3+jFIh/2fJoEU6i4e/n8muIMV0UmZ8yHN0aN5mqpZxCyIY
eEV4da55OHyeb8P5iMuwWBSVxlYTCU6NdqrF+yN2/gQIw26CaMqmKw3GyoAyGjBS
AQJTgLmZosjTHeED387keMffT6jq0mU/b0IVQIql4MtMBw8LY3jubBcJ9YnBdLXw
zgfmAK4VBi5tz0Vp6r/0gvHq9M/Q7m/8GWWLIlLFScC1LIvoh3EMW67f25Eu7zsU
Mcc+E8+jvYxDcpCXIJpvZXBt62llPtj4BQ+BVZga5K5/nLH1YmggrqZJY+VdIjn2
j5IUi8SY1P9On04MKuRz4qHRkOtrDUbf10TzUaShHdbVny7PyCfmJTU35pPmqqFm
zpOsQHDo+//iCX4s0VJ/8zZsseZpgndx+BZ07VHAsphWXi2ZuTEtBgB6GqLKzbuc
x0UkK2Fke07aWHnEQXMVAyth19wwKigROQ5W4dX+tW4sGfNIiVlKiiDEsYyshkpU
0r+WJrerWoUGZxuEQb/4eJ7ssIr0gz8cg6JejbiKIm2F5FIOxY4ynJEW8gDfVA4g
ZwIlP+gGTf5xxPr6odYL1hdtRvM7USdV9FKKO3G8jBNGEp6OdYM8P1QRvf3Vw2/u
iAEieRn+Uy/+dpPaHDUglS+838PWJXgQngxny1eafDqto8PwxzGydaJL3bgxEg4k
w8GkihDtSnakI9yU4hDf0ljZUB8DR2lQBVq1AxN/iw7zj87nZlaPq+yrLzFKkpfV
DJxrIywTh1VHNxYz6a98URDv+xQHEOha+zOCUjvucq2UP5iS9aM+I312QmlrxWIJ
LIB0As3iq9zk8iMELLJWO/5I6MFLz4dQGBsWeK6UdTOxsLGl0QBmFvwXpst7v00w
VQvtqFQFeot8rbNFNfQWCJEYaxOrOf7MkkQmu30VAbOT9/SZ4ckuK6JHOEf7doRs
wVMkTgWjem3+opVAdp63kKjWdRXM0wQAZXgy9AHsBSlvrYE3LT9v2jzddTZ2kDYa
PHK3ezRIagaS8K9R/JFqx5TPNSM6Vo/ObJRpZ97jITu+0IFQ8lHgDSrP8usTavc3
yFmmsa+2crqvQ3FrRFaotHtIampOgFEuUEwl3lU0Y/g7DVJc6gO3+z/FwYFNofaS
c4SfMByXVIjDLodGj3hXYIMZvZMPMSlIUIVJwOmp0K7C5aqkc2EO0K7sMmPfZckx
anBgO5kxJYD06bqae/4yUIMtsBtPc9V1iPtZ3Q5NN3uZWNnPCbqxkdOp1Nq4IK2P
CNf3ylE3+/NLgS84ktAloAuLgMVcWp6mLLJFMNTNQ2BGb3P6MDTWWdDjuqbHgVZZ
huFx51nRxgf3uhDbAtjt+m5p6TMEK/C9L1zovbsVEODdNVtRJWu1tFXzPz3k1xJz
VGo1bfrCyzP1hB/3NEifj225UwkvaFYwL8+sKRtDfIl2suA14L/oSg7sg73Cmhs/
vLnM2AHsvmN+p2J+MegAbfJHOQ99wYWuig+x4RjQpWMPmEVy0kv66JtVkfMeGNuu
qLIiNLm7tHM0mX55N5+Lvbgqmq0igJP8SDlO48UYtuvCQ2wli8aKvWZwxQoKPKNv
mmdWy1/3EwAvUYq64jxE+Cc5XHQR9nSMnyNYtSnS8qLZG3k0Wb/eDTiVcbsOg+PZ
5i3wlmyJat+2R3MwXXJmxK6pvPtaKCKUfVc5Sl05KmHGBMCCsEHGDsz4N7mCmfxI
t+FfdggiRqzp1Xc8e65Qer2NO2QsIUAKKu9Xl6oyQwRD2HUvvwpS7+gcXTTHhUyr
PYFZJkTCu1nnsFaaHE+DVvEuOfivwVHc8bqG1V2e+wsgRTJzktBCFseQtTL32XsQ
B1C0gjI1RYIbXBGp0CT2/2QFtNrslwmp1VqhllDBNxLozdFgz+c0/ED8LUYgAiLs
Imjzmw7DWzx/P7O2J1ZvOZRGQY4ahg6StHDkhFNrtN84IKXmTVds3b+lQgSX+po0
MnDnBp6daZz9awl1AFOurQEAnjn11wd+tJqosOIU/WiIimTAXNoMnZ55twoPb1LP
ynabMhtVHz6bCyMl4UGmc+Aas5awtVDNxqeOileieA9wvZnHrbXktQgsWqQB29kh
IDygjUmD8N/eKjJLKzEInThaX5IAqPqYuU2wSBJxtf/Zc5PQTjzvRihw08Zg5FAs
/UWbRFf8tm03p9FbLAEXSKIRqCFGLptLX/TSOqzM/y99i2dka3p91Dy7RSexlOx2
TgGJUx1qL+9nbB7xq6jL4W7dxXC2RqQ0PNNXHJc2Eg5SwxNIGDRSiQ1geE/FRBHU
7KUXP9FXcX7Xib3vBT2S0hpOtDpBEuZziHbVqyV8TDJtZ3UwOu1L2WLC8LyyP/Vy
keuPb8A1e1cbfePgioQ5UYpWEyfYoa/C/FZARFl19RU5/a4HHQ0ddRT+9ZzsZkJ3
5aDJvi8xXZPgZA3eyO7NtcZAcZ6I1XhXt/WYWSPBXUO41uMPOl2a4rhiD11AKiAt
L6DkUvEo9zFvvN2bbyXhmYR9Z/CpZ6tRzp1Vb8rkOEtTdKHPbpx7OSNOPLAwwvGe
+Ng+dRehyQV55eiCSEKg1Z+z7lhhkgL66tBwY7VQXo0bod8JcKeSvoCDVGZAHrSx
CXfBuG67MJ5ScNGe/luAZ0FXVghrn4Cp27bJdijuNY8gwF3m+NfPKSBlqHJXxeRx
g3p6601pBcfWlNNGg7hL85LaV+QolxhcoF5tyzRyxc8lNxefQTU+GFXScUrxyyKJ
UMCkRxrwIx36g1dvmGiJyfkJ+B1RlIGQTFlEbApag+PLUaWRGf6R+aPXYNQQBpSK
LvP6dN3d9yMDi29XT0tViw69CQz8iVLP3E1CpTeXl/X3QBe3wrsLExRg2E8jOmGA
yrqczx3iWeL0b0uAiDfTrtWg6VX0b6azC5iIXcQqbW/l+KLUIhosAqjN2v0JKYEq
XGN2eVXt0wDq8pHMbpZiJaDpRllTYZazLdUMg12RQU3duvxZUj4s9ASKuXy7xrYX
WJPzbi/BJFdsRwEB45uj3/CSVwZK6li7MEUtc80enIsoMXKIF2xNbkcXNRSotW2i
VwfD7+edjMnOxE6/b4WDhhnpbSodQ7ur0JGx2BShAkRhEUvD42d29XX7lXGuuJ62
Unsu5DFlEGzQMvaDSeUJuSCVE/9ZEvvYcwLAuPKw1mpSe8knWiZSVeeJ2wE6Tw3I
gbBtmv+L2IxNBy1B26MhyWZOYDNJwc5li+cunQjjbR8G5e8koz9OnEcgjeOUBL8A
f24SyowlfchHKnW/J1Wfm3AgO8a0paq6NrDU+Gxy5qM9235peyFcQMCHFr9Js/Y/
2hOBtRMf1lkYuir/1OMwC4squYZR72ket/hpNV4turHj8D7Xtd0MpTdXqRQrcTiz
ju+8sbYRP87e4VVM+x/U82T5D+amL6pd/hpXbeXyFosIj3CbcjITbI9pFzgxk4EU
A6mgxUS8sVucuPJkNbt75wWI6qDg0zGMctJ1Tz3AfZURIUjlXd32FhfoxL66EiAS
4/2/WvWKE0xeNBpztC8T9F2uLkq76FzGZny/S5hkFQgpMi+QpKrpP+GLFZC7tGxC
9NlKATpdfcTVyZauOwGXYF+PClyedMpFAP0VO8vhkUJK4mRW8u9EStlV8vkDOKeb
OFgac4tmF5lX0YWrIsRhpV3gscZjZ+V53q8yZYiMjd8gjZTIjYDNH+HEE0GxzQsM
eBFXwfnyV07uwiF0SFyEBqw/xpA/XzuRBphcHzlsHftOZlid7ml2GFjyPqR6yZNe
anOhgE08EqGr/kbwhjy4aRfngi/BDn+F+OvgM7TubBCK/E/zTpigq1fxpHdZoh/Z
LUNsnTRd+oeRVYoCb5CKcBzEcygJ2s/RwNIAyVEzAdrfT2xUKtzgEc+DKcmFmWZf
LYSjH3WfMwMtlkSkoQ0Z1sO2ruKZdKWY571uuF0cgrXOucL95kwReJ4RWKWnlvsf
XAfDsC+fSxmeVE+mrbXBJUEcJuTR9TTnqfoBe4c3BjaMDqPDmEoMhj2ZKyubbdkR
jTXWTe0/JWgHjNlQYwueRnbNAOaTnzbP7Pgg0lep5mg3eIvrEuBbDl4Rcty6pb0q
csidzUeTOJm+E1RCoaiaMFwEIE9AsJ8km6h7ZLg6mig6QeYaacr5Nbzocrl2b6+1
VOdWXbvFcWgqC2Q8jT8ea/GDsBMk0A1LgTSo5ABjZUaLOvkdbvKK8v3QB7/FtYPu
FwcB3AZvr7JTYjL7wXMtlZqPM6RBJBlgPpqKEESt2MZT5/Xm4lWm0fGSfkDgNjnT
NJnFrUk/t2Hq9jee64JCR87iIPcokvkvnheWRwhBON8fchuA6Q2S9qwpW5oSNe7g
oNlRrPQ32uOeYud1SH9d2uklyJu1Mg/hI1k/SIiSmzwlHuJUpzBEBGhUtxUPyv2a
E32p7ArFjl/3CZeyqzcyjLlekPZ6Zs4rgRyH0GoaaIYQ5p8MVtgeAkG/rN6uVUcS
9Re2KmCyEhrznWZl4r/iV1959rxhwkt9ka5iPfFl5Q4d2MzC+ICvWM51HMRuPxfX
/GdPAiOeG4YNyb5fWwCeoFb2srCif5M323MX2Nwe8nQDKJwuernCvJlsfRP8AbYt
df0LS1bErFzzUDbYZQTqYbqerof6hY3PuY+lJd8wFVX1c+WpypR/Ks9QvGWxM8+8
7RrTa1z6NorzaxD8PoHXHuFbxKmYA+2ct1x994dGkQBd+GwpUr2kBl7/EG3fa8gz
Gt6dlx+Ie7x6eRZk4J+yi8fnSr5ys178DT2Cc7hz4Cczs9mQsu0Vk8SRrcUvul0d
iD6NPSZ+vaIx9OjpYDNhlGbO3ZSJbn6dLrDvQGZngTN73lKyIXK8XIQOkmBLMknH
luAQ+nH7CPMK6UPCcQbYhAfcjkVzSB1eDwDO1gMPidMFJChkKeFeiHNgb4vZmqoS
UrrtMwlVni4JQHg1nd2NIMvnPIGVgFwcTsW/fuiM+r6rnugoC95yK1M3iNywZmeP
7p7rO3r0Hlk+fF7DxR/9l5sBYGr2Eb2Q4CwMlPwHAKiZsdeMdEW8NffvfgH1ru+R
1X5jJL7RjdrDwn/ZUNgz0NJnAl2c05TVjmjpSpSUAi/Boy/1JilfGZneCDILP1Zv
YxNMrTUi23uachjD8Ph9vlP52oO1FvZae+hcjkM/WTCA/V5u6sNjovyyeFeiDR8e
4RuOAWxEngGdMfsjBujjfx5Gu/P2taQsXuGqT279ympW9q+VEU3lp7hj/8vnFOpJ
/QWzOYRS9XpcqcWQXAg97SC+asnPactMIn52qPwZu8ETpsyXPBxR57T8kg5v/e8s
BcDGBvdC066PGxhrjvXah8655SZ1SsFkE9edgvmRptor1iLN7yfRxE10vaYSlhR/
5GIl0dZVSr+XtVNj3+yezPOG/KMuRv9FktE6tP5PSNxQ23fIxYFmmKtd5LFYvGFb
iLVWbOSdmhcxB8/GwsCb3MrheoSv1znlXXRQMwuSdTut8QAYTd0NkfnzitL07XL7
RKXwD1BNMQ2t0NCDGyoxzMpCH5sbXn+n6tJjTYvFBurPQ5pxkIkFnL7pFWI/QGQh
yEIK7BtnE6jInoy9/EIsmx1wYtyrzrb4ALMMEHtNNdL39Zrgju20WYOJnl/kq5sI
PkF6W0kCf9neqps7ZpJISqVdI6slku+9dZNQV2CmGZ9cJiluiyr3xyxUty2jJn0T
kRALRljkuw+kfXViGXYgXQ6V5gllFalrO7rQTv3YDR1LKG+rTNKrKF/1q0JjxWaL
LVQWOXH0hmygalrsl9tJgLKx5BPNuClJGeEVsndTDCQ93CoWXTqYlhATpS+5r2Jl
eLdxu7TXmougVlKVq+z5R/2G4K8mNRqQM29lzy3V+HUq7+pvWJMo4YJZ1eDSnM+V
QZiGX9Fw0oeGccwNd4ioUlbBJYHTRogOXvk5ScRbdoRCdZU7oBY9ZVqnxXN0rHUl
zOqL9oM11aZLvK9sOv9AtZ5XVyEnuKBQQwrpNlc2tjaa6qAdunAxlwmIk6dAaud5
HMdCt79cZ5RencjKHi1cJCChiXETspl6+jvKdZ7zc21/oUy3fe1/TtsaRmiQUvkn
+SGCPTIGV0yzifdSzEU9kfRvW8qfFqcNYPKqewqeTUxtJ0miz/hzQYTGJ7N0QJaT
DRS2hA9Didps2LIRKDKgWUb5iVt9JKv7lzoTE4KulI4G4pgcDr+PbIfwUWppF8ZJ
XmAKUKhSSphZD6ELtUrxBEdtD94OB/KL/N17JHmjcDm0YYPq3v6tpm8m2zRdb6O3
iNPT245FeSzH4A5x0EBxUHk8yizcstcj+PgTB20Knd9HdXwfUua0e45Ps1yiQckU
IrUcGq8xS5ui762KxWDR7fFEHA4CYtGK5EWQLmebvNb8uSAzETJS2NFsvzn1v+6f
8uXClsUNFhVOk9JK4n59EvBMk8bNrAHLS2vTkDJT5HAECzzSWgGhglpC5VwViPdv
aQVpd3goWTB4+WFxhxxyirUqUF0THReiywsRg31ltFlx22b36ARJ3usV9KF/4X+4
KSEvGFPhRvXmWLsPLViXHNPi5J8C5iERhgsRPaJfMs66Oo4tp2TzOlbwK09Otfrm
hk9x+CrWEe3ylUP/viOoRy1VM7mAbFvPx1TR9n8vqBXOVNlOrbfhpRQaQEKSMffG
2X6M0ZvL790+Aszz4nHEzUElN+7agiQ7a6FoVsqcGBpPMnfZdYPaZMPIne/n8Swk
QHKvAprgsMYcNPlrn1mjc2eaefHTwGWLNjnJRZ3i/a7Xi78qu4LDXP0b6HQyEDuz
kmqRAaFUiPKTkW2dQqzXqiDiyaDgHcqQXeT9d9N02YoJ9hfphdrAeKjf0IqQTUxX
kH9aHsScdBHBMNVIZF1ien/eIzbwG8EzhJ73DXNa7txH3pZGgMs+IgvvdVmCPg7F
5vzrakxT9XDXBBO4N7N3lhNpp7vWNxN4zdoqd6fKDCMT8aX92tV7FWKEGxbGkEv0
U5pA5WI0xSpt3r7+sgSFwYCJMtEXEc1YaEb6cAZIRyydycmikU2jfA854KKazi+a
7lNWxF5BlX+hlacXe+GEwbwpPEjiXNkR4j0UuIgLRb+Bcq9O++QFNGR/2c++wuIA
LT1sb2p3t9dej4ceCeksTNvP5NVKDmbaQ4N4W/mECexZ3GhaEdJ8tW0Au8LLIROD
K6YEuURAH6eW+E7LfzhcHij2xXzS0kyILSz8I/J9XgJlvH8+mzW8kwHYLAwsb2kk
Ktoxjpu320Lr0+onX8x4O10B9brTVPuAnA02S85y3ebp7ONIOgekhMVTULtQz1dt
kM5X8MX3h1JSETNCytPXGA19IdHX8cZ5xJCX3xPPleqysoS+SZx68ye49e2DR8uu
eRApd2zWQZZ7PpJUKfQ2qFqNkCHWCfF5/mYpThbL/ChAYy4xvz4WUYhGYXKNelQd
QCcL/IoEA4pYEtETb86o8Fa4xqH/yhTLXNAr2g0WZORM8G23oCRppWUszTf8+Wmo
ubgX15AE2Zp5GkUFiy5pkRPLYfEfN0cb6k9fQfdJDoQmVlKCqkZp3TVJ6IP/51X/
tPC0Zb0TPtSuoLrqCzmGh2vMvqWKZ/T0820/kD84mLrHpabcFlvvOcL6zLwgRFX7
f3H4GFP4RaKewd1NQLE3/JH08pczI17Wrpo+D5ULATdeCaIVyE3TfgoQf63+GAQL
9HSDHaZm7Z5xuflfeKDALxDzlSY92nm5Zd/qapjp4BThpHBn7S9VAd5FEr18N7gj
tOxRYSZGoYdKLGsEOfMsrxo/png9x4wU6J9LpLcT4sdPdLxumZA49QaJX/kebiEx
NagFKLJATwjQBkyXCs7ecJXiRK9px7UFCK0OAMq+XHvZHKv51EgG/m6NZs26UlWY
t3tC2lUB3bwd+jFX32H0BveMY1TTJdhzkCOl4q0mfyOpYHZPzrbWl+Viqe3e7oGE
sXKeNcMTEq87KRc9a9q5RSSAMHzQ9CM7dsLmJ6K98TLL0aMc75OMW6xzHHarQpzv
yzckJ2zhqOL5QYztkA3O4UZxNgD5cdeQrUd6k7r9aNaATdn0WgEPdbFvN3pjuiMc
0Q87m+jL9PYZyncUthk9U8z+Z4vWYGzWDHqZuY3sevUTEK+2BAwtOvXMkdCQcCnj
hwt1JBFH/5h/Bkx/k+sI+zE2V+eLXhQ6Kxeb6MrHPLi4R5ZgG04AFMP7RmCSLx/W
LBmdHouxLohy9EjNWvIndXfnnBGUzWsVOhh6WVRhi4P+F475aEnPJbIfpjSWgoZR
wtmSoHn6fwNuZPzydzQ703Tsw9AZ74dHL4nN9sjapvEkr8NgC9kWtpM8sS93NP4W
XXnEx3TE52rpK8mzVvF6V+/d94Pj1i3qLNqDxPZLwF3OYtEWlnxjqCCkWiG4NUPd
6i1gOL0dFT5IngwfJQIS9y4cehZwhlBYfpcwoLQv/cHoLl6n36Dp4Wr5ScuXk7Yk
7QmH1unG5nY7bLULzD8DoxWwRhgMatXtT2AaD2EEQOJEHXXHwsznnQPYdCZn4hSb
gO07/XxVeCk6ivVrLWcDHBZxoLMY1MQ7IZEnkBqSoOfg6lZuX3X4Iec1eIxu+maP
elV7weHEPZZKJTKYhfzyGVjxYtjQVrCN0QELLoleHEajq6bg6tD6iUZw37Npb3dZ
ugbOtetATQZqQF8lar8KmMGFp1deJbKZmGTOF/7dLInzF+4gr/xReL7PrEQr6CbV
VxxHY0lhlN+8c4oAYik4ewwNf84ZmZA+gH/4esDOMNkqRsDFc79QDEAKbjBzWeBO
KrlBXKbDMcsg3GP91i5pP7rgE8p6l03OQGLzTCMB/LNB8CITVvPig2Hm2/+qRgvl
EuNxf7kKf4ZhzqOcPkA11Mc3X8phEVtacSxqE8KAfYCFRqlzDrVIpv68NEeleH6E
ew0zfWK50Pok13wQRRvIQWxOh172QqBMg5fY+/ftZrvXITtBrSkZTZZpIAkroQUh
ZYEC8DJizTCZmXbE8/QbMMtVU8L7BRz0Pc+6hCckoJXrLGd6nplveRyZbL2uJn0E
+RFVLBJ8+waYKlF7m3sRdAiG5Kr/B9INPE7bT9Zga/S1h91jaajMIrLaRIG7RHBc
DMZHNGpFg/oCG4Bjid6+wk/DFWvNzeeoHUqCl0bakT0kNiZ4dls4y5RALGNa/s2P
bbNPcUPAL/HBpyEtuzpVOR3vzD237iwRf++GvUbob41WD/Y+VrroH0jsWNaUC9kV
AgpEiu9H7zgM0NQwIPwStOcv6gMqC7Fv/p6X51Zrenihse+YyjpyoGJP7sri+dMe
FRpsZSefTmuVdG/QaAjgnKFxseWLs+FhW6Sr2VAzFC3EMoLSrP4cJH1+YonivhfH
LFSkuxZ87tx7CWb2lvJJijyW/jQtwNhhV4TZ7/x2Nhdi0rVrHTxWU94xH8ktlmdq
TdUbIs0NVwgyINE5zijtBUMoLoH5+/u6v5LoFvFWDgZ0ArQKKEMrVuJx4kG4Mnvn
ADlx3OVOgwtMO4qFqdNNrf6hYwB84LLgvtRTbjFiQF4enndxjZbOeNAmXFapkBFi
qm4p7ttIWIUp4N7z09ByP70Bk5YN6Kks1RAo+XoKLSgh6ZL9mWuTVrru99xUCHyn
OeSYv1sxwftM9saYJeDSm7MRVRstdZiELbRjwIibU+gvdxMTfG+WnXdI7wH6CxWm
yU6ZinlZmTQXa8v5qz6igGRUkwI65OMnkPpD4YWK6lAliIu9RbtZ6Iv3zZO2UqL8
1Xd3Le40OdKo3AIFlsL+VLAqOoDlnwTXlE1HG+kjwU89MJEyrEBdzNidNkhBeTwu
71t7WvgU94kGepXA9nxEHBZferwnn4Z4dEQYi/7iY9dFZOxts7O1m8UAdbbg30pl
bJ1RFpBfREN9FpycS+tUEXbRDa/6HgHEr5YlT7HC8sXNETedPEEx1u1fPV5CjGNq
264xvfJwl9LCZ3U4K5zN9vG/Aam0Pxqt+wZlllD8zuQuv/idHUifg73e1p+QDKSl
wlXQBLm8Qi8fGR+G0NBwiRLFhX8U1OWF4WmlSoBuO1OykuE3HTXu/ncCCQrpwT1A
EbsA1nSik3dLjPHQirk+X0abuswmbx6XY0MlQp2aDZyELik/Sye5lUSBxTJUdOou
Dv5b3BYzAp7NZSZmwUnhzZ25YsBFRLjIXCa2V63FqykqA5gNlHdKErhWx8UCuwty
G+GT/WEtoYGzUaxQ6hCfbx+IrC2AwF5X0udVRFqJrnDWgRaqEEE4+Jz0osnRmjWZ
u62l8twMtcfFAmfHJ8Oq7wsY6e463gYflO9N12ndsGVsc1qr4syJm1lhDNiLG+3+
4vVoBaTncxcabgYryiLi2NxK/dFZ8ZNLVOdTuVsEhaA0+3DFKdKFOTpRpEfNNeWI
MjLlmuM6grfU0U78q/ekqNQ2SGrMvY17WhXo8DrO4mk0lwaAtZaNjNrXELBW7YUP
7YnHB9P3/Mv00WfIB6NMb4ipkZ5nrB4rJIPTgJ0A7QkyGu++4kNh+37dXJfV4zrr
Ul8Ih3EgruUI7XKAcj0h1+tobPpJlaAIIdwa8Zwvm1bxour6DCzHVVoYZFdD5+Nu
HrDZp9a9IrtlR6pswHZmM1QNt4e6E4AnY1gu/q4xFxqDxpyQ7Ic7ZUOg9GISoKve
Nlta4jcSrNna9o/69WQxEUy8Ni6Q4+lsqZ8FnokETEEb7qiBsRGVEjP9NSEszbaq
XIb3bWAFcrKVrde2GSKflu3RIiAMRbIJo/KL8YKk11pLdZdM/A+qEzPPqsd3iW+l
fNjau9J0waVJNJbEW5ejU/1dQ9YEt8SFbPBOhhg4xvsbaH95Hu7sqFWKpdrpyrmy
hp3IewaJESBN7e4Cp7TWzUcBzhoq5EhBk7z89qdRK30HZpIR+61NMN7uVfAtDBf7
N65llDL2t38UDMA0tdKrEswWXMXBOra8durjGAcS2DC+9isPUitXjMJPTt1B80Sk
DLHBuf4/QNPmGZ/v6Zpm6k7vXa1dGKBZGFggspWJoSxKhS7M9bXsycvbIjzh2G9F
8UdqwHsxUeRhso/wc38f98dKPXUYj4oDgGdhlDJYrzUSgp1xKsOaSdhniyD+XJ1q
pVJ/LalgntuYJYuRttIIo4NtSlFwxZT24brnhBG2Ofai2vvmd8NfItlQV4kDqEjm
QBZ7zYpIrkQY/bDv77U0hyzw8UajsWxAns4rfBZgseXu471t2e7Pux2MaTomQj5O
iqgZjbCvMv/QtH2ok+YWJK20stA3sUCn7xSOvuAoi8F5FqOEqoKPyFV+AjgqezwE
eXNonQD7gMm2PL0KGAWpcV+cZcgo9t0sIhEgVfQvMr4m1JkfmNF9VQSZBjRBkyde
Bo2LkWxqT1q6APfHGhCnK2IWZ9JsHr+LSAPfYv0CXnKjGF4aOnsm7IVzefjtqzJa
5WA5XmBkX6IehQcTRRvARXZ9lQ93dnBZtkdBrH16dUoXjlpwPO8rOCrD8y81r0Qe
+0x1NKTxSF5U3JJJdmeyTfXr3ZqEImyYfhMpKHrHXn8K4bnhfMVGwCHFipxlX8cJ
T2cC8lgjtihMd8Z6pc6oDnKIV2zDOqG0wD5U0tRIiBDCVxqMw4HvgAH83jifAkzI
Cd1OVoUnUZbU/yq9mxGOf1XtFkstjDmxmCsce+eJbR7t1qFbnuePTt4X0M7p7k8w
b8Hs+yNLJBgNj9jWvE56/HeS85WDoQNeY6W3IweRLpT4vPCCG3QiXFvKLyGHvCFJ
uzwY66dRtIc6Q+QvbbqgoTrY7Rrg19JKaDqtNN02rgXv0tYiMwFaZXlJYWJgKxqe
h5dxge1YJ9jWRx/XY31KM+dAfQpnqYfcSGeRmVj1fSkfk3FWeTpFNUHeSbBCH5UX
1H0xoBdzn8CYOjx9LAhHYDpGXuy7ubaUMy39tVsbhR3Xjel8WpZ7xvjlp+1YppY7
KCH/S9dobccwSTjMXlL4IdmgHGAiq+ONiAquykXzb53GXzYXO9anADup+IPPh1BM
9+FFRSWK414aI6bx762KjkVX4wmKRcw8QZ6YQ+UP2oqwfJx3XAAzoJ3W1P1UcOAh
xF0jOhis6RlbLD8npc7R2E28C7WvEJaOoEH6SjM4UAG7HGR3K1qPf+e6fD5Uiaug
Yzltzu13xvOG7SMl3HeJOuiyheH+8WSylGJ72RtMPI6XgKTvcN4pjRXh4/WHfquM
DYOrDT1xuJdePk5on52m1pitPvQxcBC18WbWzfTDWZGyK/HY3Ub3CvM1+THqUI/B
f9nl+TzABjh9FZg+DG/jxTiG+VgtBjDrVCnAfGxmYfnWQ4acED+Ut4lJjhgC7LXy
rTlR4u5KSGwmRgVchqYzhoKFcHiw5MtmpcsFh2KFIq0f0FobuB/d++7sfl/xsP4s
IRkduuDxk5anhrz5fwUvw4w78+loB5xXlyU9xdo7Dr5TzKxYpUNIHRfZtL7oh5PW
8DL+3dhIOacBNpIwr9QQns15Na9zDtFLlZ6q3mdmMg/8RbRK2GvV5AUGeXu48ECp
Aw0jZB8DVwIcKgrhE6MvWe2dwC99lLHgaq71Rr04CY6FSwQdmmqQVscAbKPf9Kan
Y/K4rALBW7MpQy4bPgCV5Q3GdmsSZ4lojwBK3jR4nWZX/T+B6oZLcqm/5jpEKdk4
ayKiAWo5hOOVILBe6YDBAAmplCamQxUJCZVbkSHihvG1Xetz5MvftAUELzOtKjhu
Seq4fcAEN1rHBuVsnWurUfP472MBiv8qW2hRt3dZK28HGlbd1/uocZ4/KFLn1M9F
CST5IziToxx/lED+OtTYBQvWw1AFCwyjRNUgjpPDVwG/RFnGI3r8vWRns+hwQ1tj
pHgHx6BlzLcZ/hALfRb4cKb7JeJryTJDsatT+wPyxHlu+YXRe+KejjqumDAwrKPi
b1fszGu405xUFcW/MskLqxSE804tIVPxK34zRUYuw1BiLXYXHFXjY+gxdCyrh+wa
4B2pD0G/kFw/lXN8FG7OP4lZtw3YfjHOwsQImeSaqXS1IaOKwH6YTbBFAe0j63Xe
fA9MdJtptXZN9BOu+P9kd1LhXSbF8WtAdFXzZk1fIDXRFlo+Iqs2Wt5ToaeQftTO
pDEJjFTjw+XUINwAGNiq2j5uQsQ+y1foHBUHswE+7z1H80yUw8yz3SkPNOYoXD8f
rlNn9fGaNhiaN+ixiD80bWGn+TWI9JU8jqxvddxrgu6fixzXHFBgTvKcrsVfVsDR
NVg0jHExaBA1D/I++9FUCgVTAl/w8Z3M16/1FoqQMv8OuiqgDB3EIcQYzS8nQw+g
8/YE35pb+IAmP250QeML0gQw527L7WHSFnf6pNnlcBk2G7l12umclem116KSPIOx
GqehIvbp3O3QECZmyE0cXpAGkPWG9kbiSkvnfnCxAre2jsbHvDEhXisk5AzCvC+4
wcj2v7M2PgaQ4AJ77MZ9uGRwz0GVg2ki2d8Or5j8yD/T0GmrbVXs3RhXsIFHwdgz
x+9rhzIgQ0Ipyl0ikVUrwgRrBn//5gfUzbbnhOmBbVlFuWsSHZiuRtZ9suYc1P+t
Jvyg9IXdlV16e8na3HnOA/cUFxNtNWMMDF98anCHUyFQnxBPZJN59p+cv7cxUmgV
LrOO61zJz+salmnMN6AFPZwE4im2gLA7/GXFgMfJh8kx1q/rDAqyPX6nFhkYzyrH
9z7t29kCAxFewLszsyKH/UoeoVrS2HfjPcdYdK6Z0ilHGls6SS1eX5dkmxj8Lxry
CdI2R20YW4yCIHJ4VvBFKP8XwybM9P0yIojboxaoTrV+96NHcNJQ62o8HYlL9R9B
ScH8CAIMZGogvCsYnW83RfYgiz77M4fqMgpTjCBgKsTui5jQEL+9gXY1bjzeXsZg
v318Z9riKXAv+s7AOToweA8V4YFVCuw0QGd3i+U+Y5NwZadCLCtV4sCpuBglNVMT
MvdUTGcFKP3wGG1h6cR5GtFuLRfd85F9Q9j6x9hEgWlr3heiV6dcUYZ2h65YGLco
jOfvkk8x/XPOHJuLESeGYFebEQEB2W6fAsIopJgj4XbMf2BKxKVXzKhnmhH+dexZ
2Ft/oSQcyJptidbkra4PTGdgoqth1PNEaItdTUHIdHWpmfMZx9JoIZLpHS7JHuwC
k29AvVKAij4mfLJlcL6smlM/kcpG+KR2goXZcwY8ORg9dyZJyW+v4a6cKchMlI+H
SudofFlUwUS+OR88/8/NQAJVaTtc+d5dUMboXKJ42Nh7eeS8Z3eJdvvWX503CPUc
1IydS9Knrzan6wtMfo4gSs1xrWoxteCr/q8awe3ntlNbfDaYfMUvFwmxFz6INmNZ
L6qWf0mD1scXIYJGQP3e9NC8omU2Hnm/Uf3dx82vzTpOPki/qeyD2Kwtru451H8g
tACsOUKGX2nCjBSgLtnQ0eTBVxV+FUY688yai+FMHVeIOoTHa/EbN4pFGcx96toX
bE5XzXBw+h2EfFy5URrBnSrzBMtZh1Offyhm4md7anYF27rh5kN0Hgn9/ED7C9yB
ra0Pmx6U0zpga+E66+LTRTSGJl0Cm3U2uUVz2rU3yCCsNyA281DH5gpXP84ziy3X
PZ4Mg6NGI5YSWtnjB4X6PU+MQ0e5AThCasnHwGC8XdccB7en5zUwJZCUx+BeQZ8n
0KUNJPr/3T7ytNtIo8Te2SJ5dfLn+BCYg0RNMg9L+sdou+YUMzF02JTD2z/KSZ44
XGCjdePrLyQnGDW1b1ku8l0966D3O9ulIBd4uOsabzUfKswLiU0prMhfCOqnshr9
IbDfWGuFJ4IZSfiFc/YA1hbt1mxFSsT3FOi8DcIeTf2fHxXLYMRtPIU0T60sb+BX
72TEi6zbyd4wyodFRhWtzYygaQJHzEpJMhdJlpEUXWWYNVi7ku9gvLXx1sI6xRXS
iFYnN3Fv6n8e6cgXMfkvY+xkR58yusxSSpTARbE0mva9Kr+j/n4Yu+tBvVNxFOsY
zbnUp8RMGH1hZsD5p442kux3x8oDwhhHuh1YHnLXFHmrRwABo1DaZ2arFLIHfDa1
S1q93GmnS+dVuX6BbKBlju198YjYqP6L/BbC2AZDEvwUUAiXHnqpYxrc9WMZjn76
KyIlbsv+zyEwxCHyG47s+a7jfgyhyOtgJnOsrdpc8Yy2aKogat8WROi8l/sfdJ5g
iku8AtWznHLKs6Del9RlPY0H4qSmbgQYGaZA0+ayHfl43MeNY3cXyW2j5rQFaDY1
zFhXpf+azZTb3lE1QArthPXmEIVkSeVRt0CLYz7Bp6T9yDpUEmst6qikxdY1IUPs
94gCrrWBurWSVCHjwyD2vSfGoK9UFdLbRKrHME9wOrRonapm2uTnPNZvJ+aGqk1l
K16aiU2t5zCfVgB1L+yVbGafa/kRgbcF6vRC5XLGx/mZADR1vlKF7gwmD0vds7lz
I3E5ypEcezinOj+WfsCmJ2cB9CXwMh7Om+lNX1BHOLeGQo2GZUBrRSnjpnn4uWo2
JfASLQEiKgQZTYiP1VAyGJ8eyUT3UrqCSkcDg29R1niV/nD++IxwTq6N8O/YzCIS
cUVTkvrt20i6dlatdJis/o7e/WZlw/ZDzBeAbtHgCJ3TH+BvLZSsX8IEPNZem/sk
St/+Cd77f7bwzLW5SiTKWJ95eNu7Z+OKjhM305g9Sg/qYr9PcGwiumdOhaBmjBj+
B025zgpRcZK2+yGo4IGiObGRUzP9qO6UaehXfCw58aWqHyLXOxRr3wcZGJIRXqAC
3apRs2oAe/zR6464U6QxXmzHnNEq5Nw1G76ISNehVD90sw5CDxTIE8yOMlDUI6pg
LC31VN1OWp9e67+pxDfVNwqUYBHG1snhkonuGxBK4U7IsBGtdIiBiJpBjNrEK2Sf
h71c9crcFie1RbbDnz778JIOsjiUUMPrF0eKFcv4V6zvCmGgNFMWymna3NFR3471
yf3Bv+wqqD/4RIOvpVW6/IIKVFh6SD2SMaHbhMVBrBnN7nc7T0A/Pw80ydDTnNrw
1/Fc6JVWHcYfpbROg8dcubHE8mUNGnQtyKgAdxGWrBMsbaSJezGwLSTkFUR/d1El
RJ50HdwYVr73UezcNR4msrBwk8t2l9Hh3PEbgR/HJJQFBAotYXFTbYnhwPfJqVF4
oaE/ryzkmp7+ZnR1sfnZYk0p/xj5C3HaOafNLcYEWtjkq+J08/Z5t56r1XZ5CJn5
OAIkHtKn5Bh646Z+zp8kUC9FtPzoeCaepPFv0RxxciYPz6omYJZSMk8z/BL55p8d
k/LNs3WQCpdcFlh8gtMehqSlBeIYIjQKyS1jbvo4gp6eiDSOQqcoyUkTwik8MIlq
uWxBk+VcwattGaRipO4sAQ62lpD9a8UPyz1X5TZHh/zYO0oMvHrgJWnyfvAD4eaR
Iisi1CBwoV4jq+UKzMum5VA61alpotilli6HW6J6/eOp5PCRht2kAqkmhiKFXvKs
ZJdk/aN/sdA9TTPeKIUv8FvGplZ+y5FYHweQX1EleKyANaXz9cE8xemlk6pec316
HLDsID8L3ImpvGuLeNcHaBHDLv/2UqcqRWumUDlVg5fwWbflWy6sNxjDkp9SPlp8
JY4LdhzTf2Jq4VtEe5ZHtMW2EmkD8I7AujRlxPd2u6/EWpcnYjGpPfNPLhqdtQOu
B/Ob/k3Rp9Pq7uGMSpkKhyY4LGGjN0KlWrkBmBH0ZJAK3kFK+UC11eDxHxhdu8sG
IidcJOic6gwGZ+scgaDKLa5J9KrT/qMCYQoeGWiu5s7p75gaBQTGXg4QQVtA6VYj
la93qRlL4zBk/Mm4Umxa5eX9F1L0yZ+UIG1TLUzkrFG2i79lc7KOFIZO3yYruZRF
HLeCs6n+6bj4RofQbzxH/w75e75072Chl369/tgJQmqF18NeSoPwefGoBspz4Od7
NUT2tScvBX9BzuVF5SbNV56iHlLnlAfCq63oERPnFrUZTv7gFfprbmAsOZWvmnSV
G4dEtLYAYzR/l6Kq1/d54tn/bKuUq5IvwnzpYRkj15gfAd5ZgnxuFkk2DhWnWDbV
CAF9qOd/eKvGWpPi284BBbXrA4ptFwZrXOICjdxEm0O4j1rpsTkV/qF/+5aMimBa
QvbABElVuX1nqtur4M3+THbP1PggZMWScUnACuwWS8jLxAyTWltJ+TXXKN6D5V/5
3TRI82c54yz1w4mSTfGe302p5M6B4aw1E1gqLGNmyVYAivFSoiEXY3vgqvjlPpoV
PB5HkNK8wsLcDc//rFL3f/R4da/c7Y+sBXY69s82wkeFGoGkmwJjAxOtRiv+ni3E
7JMCjbVkvclsX5SMZm0b7WYOCeOj8Mc5rk2sgZHsm1AXBL0Bwl+6Snke2zHjQYG/
/agiWYo29ooAWJ+90umLl1rLJ6IspU7moeXtIjHOkIwojbevgOuiZ97QbXrmyjdm
egch/60pj5LcdPHbQv5Zj+PwikzGCbpOhdbL1rvqlzDfVOUooqu0lFCRmSbCE5TB
igpRwtlRe/T6aWwFrgrq0A3s98iNiD/7Dk+eZsPdxNVokeEtgc3S3sXTRxZZyqF4
h9hUlpdEqh6SAuUdrVvwKl829OjMH8H4bh2VcaYQDz7drreFG76Zr9v1Ionr6FEa
JEAROO1SdbqEbkMOX41P8hOqIArfHDePVX+Aq4K2FIk9leUFnncdvhfM/gTuxiV4
jpIZx2VoPoYulxsndO3Can8WqhTV9njU6uCFoEBdNz14O30O1c0q1jtgk1EBL2Cq
goieZX21QtLkQUn0uawQvxnX8HVkdCP4X5xnXnEIHTstuXjF4SClb3P3tb2++tlV
aEdG0Ct9OC/v1qsiacD1P3S1MBnRgfOhPYMFCI/cFrQh8WN9cBc6sI09jbTW3HZz
w2fSr7rlYoTo9vDxWprKVLM0p62L6BrlX9nnqu5dTuAOtOUz5iOLDuKJuxNl9IuZ
GEZNbw/5mqFOZiZGNAkXVkd6TCxrS7hL4p9FQ0XJeR3XCCIEL8XZ0/DiSsGFZgQG
WYgDTb3CctvzBgQhMmqpPng7WUPGl7A+SYwkjV2AjbO1ry8YWwFrPXjIoG5aeUrZ
yRMrmkuESZRM8v2+ZAaMvDzjoNK25gmPpAHldF+gtWJ6eZHeHz0Kg3q9uAjUVwol
UzUHltf7bIcUGrKE4qPiCEtmOIEKCbVhFxfmSnF/dTAE4s2yT62W8uFzGl4WQuLh
by3umneeO8+6828zqpk+iREBKdeeysKOdFaXWIJrr8BXztMUW1fJ6iq1AgLdeuA7
yssV1xiZQJxm+CCEgeCJgNO/AcUFhqKYh0kXz4vKjeQJHLFoMAtRivQ/NBgTmM+F
Zmar+cDGX+cwrY46MbxWcU59wD/KjdFx59/xdagOlVtiAKQv4rWjVe5v3O4mWw/C
q7EsGYn66xN2AOfVkyWqVNF4Bwrvx16cj4X4z6ByThsO97hmUfT2Hes4yKuuzshV
ZkAY36Epo0vKnF63tuveruYnZGvYeTyNqhjcmCLF69S+OxvD+1pi20g348/8Qceu
VeEsV/pIiJmMAHCsq/hOkWkfB/DybfyDNKZptK32WiLljHJ/lgRDMRbFAJ7xSYQ+
oHbNRvyxbXdtRp5aI/EQvzDd1fQBoSz5zKcrUHkScT8qeHUtRWw6+c6NuNEu2RWR
jGzjNNyLbD4/ymcN3+TY6VYTLXIOY8p4EgHF4BDqj11zLmpJyyx43s8mJ3PeK9u4
z8z4frqvoV0WY8yUeMGuUoEGtUkdIaC1NP60BZTuoIt1NrRhkOfCnvFKqvwZvy8R
ii9WyX/09ADnYCuAfKMgIiZ1gs2/VikvBOMiWvzC0wLlFss625+jJdAPW9265iJ6
gmK7xc0Z2dtt1IrtGPomL/BkDECkfPlni+cBZqzRd8yHsWuTK7BsEk6aL/6PzODA
XdD/M31PvpbcMAZIMazxlrh0+K+hCnLPMOEJdz4ffJOViHYFkWohbGZfHC24T0th
sx0axt6FGKZfkk1qhhuuCFOYm7exztSWSLb25fePsj9TZjDqV9fHV0D0rnUrsTfv
RcFE0uOJzq8PcPGxtZHrMXyIxl+itwID8Nt1C1pGTX+qQyojzJXPljqxz4F4I5Oq
ACGAm9gnUxkm41jZFxdrwBwQcpH6xyOe9SeWbiKl7t6v5RQK21yBYAZGSqIAT4tw
EIb7tC+A9UVMCufmKXVS9NKDoGGIx2F+ZN7lrX09+/IRUH4o6OKV5hBvuuZbXxh/
lxf5VGiCIdldZ3YaROPaMEpWZC2GnEWogzC6/LkWcTm76p2+2tgsGV7nyXpc9dL8
5JcUPGGGUgFNTdTFpviaR3cNGqMsmEI2dkf76d8h/Ze2SwQadkY0DQQpC//p24et
ZHguAjXv0BIgKkMFOfARiXNrjLvqkEiUUDRtvssC5Ua3jAByd7NvREA686NuyW2O
0AjrvDo6xCg4z3A8hGLWqDEYpnOLe4ziKrze8ZipDCUWtktDyh4Nx/gR19RJ5blx
LcAM7miNGYS/ng0Urtxgjg2CJZ1q6854Crub9Q6Ee5MxQqnz8maC+xTNlSSw5cSx
u2OGH8kb+T69ejFkCWlD0jdEWqsSmqCmQPCoO6TJwWuCSdWctk6txROJq7wlPLwl
JFTlvuIi3tpXhW9l51rQszuyhEqhPrXa0Vvd+TK7wAsU59TjsE/yCipyEvGN1xEk
Iy4U5pJ8SlPA0QaeqeTnzrmmSazFyiSOuyJImimYPDRyJQoSryTUs9SyVk2a9HPP
AXn20F/npgp49R4GRj5B3vKz/UHdqZMjgAsCxAnR6jhp23PM1kC3dKJL0hn6yjyf
MtwKxmJwTu3wuFY+Og64RWFc+pUjGBYF2aC8EpWWNiBb40uTtlDvW9oHUZWH/WG+
auqey4wl8qLDw4DLP6VHbUsEIoG2kd+2KwKD97sQI0N+5XcgxMwQBD3OLsofcfAX
i5aLKZ7gADNFnnkQ+0uL/nsBSm5lh1UwBaO5Wmot9f2EEuLRnjynAT39HZCU+7I6
ZTT5NxdirLHu3TOzOEYQDCJwsfPUOV/6vZqm84oFJe/tqU1tux1v3lsu+DOxRzVg
VtS1BRYNmKK/txIMnBthbB/SdFHWi9DpXKEJ3Xs9LMp/eyVY5F2568O5HCto/PD2
pyG2JEgPvS/ApY1cInys8zaIlnu0luzZ8hXNLu4LiXpztCiinWmMkw1JeLSgS3xf
a+ga9/J+q0sUEzxhoNHLs4PxaE02LSd48vl7UmkcKjVJfmMDe86PQ1J/IZYZP1kc
UJCYZa471ZtqPkHIdEqso5buqcEk7mSEeQsxdKtkiZXbnvq8IEzWITTVe2YesB+X
CLvfK/PWLHi25keHNQYaqGUNdkqyBcRbdQ63qisUTFzsDdfbdI0giwRnk27cObXE
Heuk+W1Wi/C9+zF3VTstYUh8QU6pPNgmWStM9nl6fNEU7IgOpyBHJlQL5TWWQ3G/
H3z2vfkuTAXb8Qdspm0y7eLm5JhYjZCsN/YVl1YPI5hjEJrMqXZFr4mhfoPbMwtd
X63oBrnpemsRN2yRFygW0hbhCvnF1xoPDoE97sahoxKIHced07gnAhxttRuiWHBR
uRdhsY+oIFuZn7iZCtox+/hG1kXHgFzW2Gemku085EHGObMX3JoY8vnarq33NAQJ
NNQowz9NMwduHQ9MW+aJlgAK1qFiBHMO/wTdtOfAppFABRrtIAdpK2oE53Tye3zY
255I2eAB6eEzVHe432ETe0wBnhs8K/yTAnWQ6uTksygXouvdQmOr0ZtFWLRpkf5H
zs9Qx9/sOUNvoTMm2sqTS9HSa+Q8xusY20nAz2GHNCiOo2CC1zPNNiHxLwv29IAV
zmjWsr5dMposiMuWSOIpvbFfJT5pvV6v7XmyuRrGj5NH/UV1vT7b3FUzSDu9CMiL
Ns32ys3YSVBYNdHEESfU5f0tfVYjAVZkXQD3+jZB5wpqD7kyRfINjrTr3Dy872Nw
cEgTt5Qq+YN0ONZURZHjJYX0MucR5vQD8m2JbpWY0i6gNf054yt3dsgjqFpQ6Jj5
buu0JjSj89A9u3IIBQkjOOg6NUpzMdhQXRJux1vliC1kxNAB0At2vtofCtviLi8B
xQBrgqnRy9AoHW3oFUXLgJ/otx1X5D3eppzxF0nEPF/MyRVC48mLCjaRhZ80Lqx5
oaQB5R3DpYcEcnWCjsczKjy6Bz9saT0DRPV/MpzOxn4jq7KKmyYbrM3KByMMsw90
VDw1i0BH83WXuMnaraUm94I+N/CO0m/sMuVUN3odJgWW0g3vjUDP+Oek7V6G3h6L
4OxA7Rv4ngKfDJP/VbMYjGWT1hOmbFQUkUXtbGMPIqq6LTb16F425fZkFa0bL6wM
IgYeaWeFwPEzdertQqYZkpnRtZi4zyQ499ndjhTwWGWpD0N9OocqiO9IMIARm55k
jglu//G/+lnGnoAWjQUJe0QTW8vJ066Qy3aIil4I4nSdfozQuXc467IzGP9SMxFw
0OrsC4t3Le1rVb/cBnonwFU2+ivZor15d3AoDlBcoLeyooDzWj/GJskosZ0WNWrO
m2xGDqlS4wQH6BOaAv+rue1744RTE9/DeBFAeezsYPaDNg6Y3A8fBqZxniXLhtm4
lzq19UghjFt4UwNEBUvBx/54UtFivjgv6HCy2AxXMMAMwA6lhLcuLp0aszhMnOem
Xopndt3X7XC1c14K0i2JVEf4zPWS7tFnsr8Fy4HYxqHWqY8/xtqfKCQCf7XOTR1r
/cW+psMAohZJOISv5QahVzYI/M9AbdlsEI92AkBriemxI8nsC+cW6Rab5dOMZDOG
wyAt5qFyd9+eOkMZntnm2B90LRWVyVz/K4yZO7QQtQw5vvTeu7z+EyJR3d6adIts
LDQ9GPz+iyDhUPmkGTRaINbJ0pioj6f+3VDcBlzzaN+z93nCxDvq/GvRz9rs6Rqg
CcW3fhvTnbU3eIL7SB/JUulLScsDgUCi+h1YjX03/6hHODvQ5r1o2LfLN0rJTSvd
DEFvUWus4GUcUoiOiz3O5DLS0LK4qKI8rJA9f7bUDmNyhbB5BaKlqS12LT5OeWHK
iJdFo+BpS+g8aexB+TafJhw9mqfuv5Mi6GIC9gW7NT1jJ7pCTrn/UXAxRuBgzXap
HWGyRif0GRYGITcyxcXED5gx7qk6wIB0Qt97GC4m6U+pQOTmaQDn5tLp+NjQDW3x
lNmJ8iINSKmuNBF1IgOMixIDKgBA0sM09Se9ju1Zz3r/ptyv5HC5H2Ib5hnKpdSC
DRI0RNGdj5X5AzbmRp/VRuJXU7XNkYTfpOhF4iWBLleY0vma7hSPdhrZFtvMIO8j
dbWUF6vp98znzgK1WBvCMdWHOvNwt/rrsFmBPhf+b7QeK2gGAnIfRQJOZDEJ2yol
auqS3rZAigWx9XYsAkJWnHP2ZY7DseCYX0s12G76FBUfVVEybeiHpIXv8wTEmZfJ
gTi99Rapwrt/DUQrV7a1AJSYSjNmOPhsCLXFyCqvX0DgbSYW3qr4QaUscZaZ3uj4
nnMT8CUVYU7Oe337Q9QRQkKvriZFRNF632cLqa0VoNgsyMPOUWu+/wM3XTNXEKlD
f3bfZYk/7Xh4r5tD9u0iairWlCwYaXYABjyPjXLR2QpmwBq/Nx1sId0+Utf93Lcx
2xJ8EnAQ3948RIEaI2LMhcX/zraW3rAglrxZhwKK5VrHd5GNtq3ARG4/9N6P9aZh
XuUnaBIVExRar8nXYz4tilg2DP27sTsuIAfT061JyDie7o6TGrbEJpx2TAWU95lp
zHakOi6BU2ldEuykRMS8y+fhY+OUlQi01n3qxkj8Q/7xmBNBCYS/m4CWiPtCyo3y
skBX2jLh5MQtmre3vrCJvJppAKhgwnsf16rUYqvaLnjouN67pC//0sW4qPbMdq+r
l4hcQst8SDUCQaQZpHB/ue9xHVhkaEMPZXazRUDjJkkG7Wt0UexWPk0/oqeaEu22
4SZEyNnUOXLRMzdKURFstQJ3Ubkrhv85Gu50LhRVA4fkOEiR+vdS2bmgRM54gbsU
nRtoRs/G5CRq5Nw/p2gLPTq9p8Bi9unP/ppIV4HnuVUpTx+H3wd8LimMNU1PStL7
tQ6ka7UIUsKb90zxUN4Xm7N5qiFKRhq7KaI3rqwDyIu/IX/PbI9gSu5oxBlckEBg
EdaFcNw7ngfII4KSTnnv1OTdlfPB+bJkpnfaJeZT6bdDeZ0ima6BnYyGAREbAJLE
QfYvNI3zQ0IPvlSXz/GxZHAzyITsVVdqu/Dc7tZRE+VAtga8O1whA+Yy8YvNPW/9
BWmmJ9UrtiDR7HE9ScCetQZ0sO3ND9404yqEDUetsT1s1+kHkXshrezz0GQMpn78
uftb4tW5dx5URVuI0JbjXgRz5uR2d98i/8wPgRjUFwokzzYnGGqfNCWh/BlSsx/1
22Wk2sv8Vz/lTFWUG+QLfR7IVz2Tmf2Cpr9YR2BFmPbo1clkuoPmX1Zgwb9zxoyz
Ff+bmQyJMELO2RBE2Nqffh6ZM97BDbF1oZbN3W9gH1RIMEzS4L0c3esf5o7vDtHd
q33hpk3r5mWliCUKOiig1rIkQI0nOV6QuoJ7/aWhlUnAUgzKNXEdEFgFxPgSpkz3
wzhQcRWODobQRdmyOr3Per1kcYjQifOaDXZWB01i/N2r1enMcoeMPcTRBigRilBS
FH21wFAxh0gQAslrVw8HrGMAi9mDpFZMiJOqH5CIW5PfU1EHLQ5rU09RWZ+bY9st
HJDYAD1iplW1a6ew6pNxpG1RUdGA92AjqTv5Hm/bXQkd7H1AUlKhsKT6jSnUWQCn
gxxu7CLsa/0rmig9QpVTrnBTOvNWio+bgmCEc9IVNo/+hFXuUYflVaTFTOlvsD0+
bgiuo0xeU+abHHEK4sFmRZfV3m8KAFfDqTZ+Zvpik5JIhlZ+6L6cz1PnvwKUbpuL
XTG1EcwNpaviuZSB5VNH32H1d2thTwqKACMzP/PH5OC9RIGFSuMrJ6kmQ2E6NgEQ
BoHeexPwF6lx0kYKVbnGlYPR9so6FL/et38AowCP9iFKBPpfR1zcLslpIkeHw+dg
kmUrdIEeofGkMFqHSUxzlCVfm1YynBMMroP8N1W+nnuL2/AbI8aFWpKt0s4LCvvN
iHqKMOJLZKkDlYLlPDXlHoyDzvQ8M6PglSRk8VMhTeK3g42OTcZx/VmeI2FdEcT8
OHfq28ofabfe4bu/iifOAZKm8DBiUtwTyYxb6QqIN8BsM845PB7AOPGGGIXFT0at
LQ9OjBsSvitUQkAXb0VPcDEAPSG/GFbwppJu8uRPvrd2iIOQJYt2MIt+DAdwz/oo
aHpsGM75iCM7xh/I++ojhGqq5TjgMFFM8atBCKHJsaLmV58NcrBedFZhJhrntV01
9xTIU8pjPNK8WiidMExXDgHPw9PMDAVHvDd9u+4G3/2fExfPkODuGUhHgiTmtJQT
2lEAYKpF5iX7j8/4JDWarQiuoz3YHYqYcsRQtffEbxpX4C8kpz+CBOtvp6ceaTjB
2CEy+NgB+Yoergz/OBgJq4cYa/fZBagBEb0ZWAO1acHb+WA572kxCu4vSJoRjEDt
AbWJ8ZIYWVuo/GF6evj4bP5ne5shcFXDX5ShsL5zeNTSqXqIKL3BSc2S4fzhHKpn
UwGuJY1xQyfmQXRCoJTLNa2mcL/owa1TEQV19z7wBN9NhRp8SWzTDGHCGGb5l7lR
X4i9DLJO9ys2A5MgkJHVdSd4P7ZFUESako+/BkKSON43UsMk0iB+V953i4OM5RRk
HxUAjJKDaeb1juFdh0CthcbSxjgZahrXY71YwMFi5hZm1LZER2dX6sDEXD+R5gD/
7hz3UwxRVRQKR90JazalrXE47xUrlyg0TCE47EzKLIjkZMTYUqQRsxlcSRUCl5dO
mqSFmMWOUO5F+PFki9pp/6yL0cF7tEbY2P+4eRAbImYXtUIF07F6KFrNoSw9VvB+
u0drd+siEMxSYhOfDLQ9AAfbCOxi/xaIYmiv7MGMwUmGsq+MovoorpwansZhlz34
UerUdnIKc/EaH/2eau35w3eeGWwlupMHfieaBBgSIYPIw7gT4ZhgTF246XyfSOnp
cskbZfPdeoay1dPm2p2SpaRLRERRRn+hY9OVlrwxf1nncJDcVI2D8KVof+jc5zIo
tsV6v8F7o7ueUMjgHsKehXoB9UhjISCLEQLQiC1yI4UTy8VN2D95Jy66j4QfkSjN
AFPt106oOMwP0Uze8rXzDeOruCn3XNatdxW1A+k/vfCnXj1U6CwUzndEL46r6KQV
bnTMvgQBEwkz1C/sUtXckeNQXnZxEcnvsYn1JUOGFu75kWwQkl6VBJRpCq0IBdPq
20YOp3OuGLsQjxPfcGnZ1cjNzmFPhkkfWYC+Lem0/SQIrZiSp8/ItsVZEaci3vWB
9HBrUSRdlYzft+r3Ds4ZlcDzJ7vKQu6n0Ui+hI7ssfV8TmHKZZS/nSAiz0Hs0lQ3
Oa1agOVlbtqVwaXD2H59rmTo03hkrPNW8pN4ECtjM/v02OHY8aY1+qK4Y9d1KuHg
ZtZkHuoL4tmRcr1orvKeeTJPkVuoECt8KAtY/BjtVDHboxg4mOAbsPuaUj5lmTZm
wiRuGB+uA4GJf9riNlnh1mZgrX76zsujgNZylLPnqvnyHb9Klt/3QutnEzdSXxjA
7S1KlXULQfz0O9meJhbJT/Gi3KAc4iHxavqOxSX3tynKFiN+QPv8iFgqMfp2cWHV
YgYK2ecZPIyYkEMaatJzz9mCkEK42t8ig4rwQDcFOdLxLOBIA14KMa5geN2eR9bp
M3Mfczxp0JpFhPpcFzQfpCDSpe17duGKiaxruCJFMRpNwlCmO4ez6MLC9khEAY4S
klKqQ4u0oXnu6mR3MasxF54TN9JZCi+nmzsLdm8jSGEi3htnZ6GvpgAzxEJq1SOB
Zdev02rIk8rM63ogWDZRSwnpIuG+zu6KyfSUumL/p0UzuvlyOT9n1IdC7AuP8h44
wMnORC7Wc2I8ugt6kDzI3QpHleEUYVjH8F2NTwVjMZ4tvywhTFKmvJr3JnlR6lzm
wk9O8ySEIx3h5bWxzqLxdAsijP3CdQ+8R5N6a+24Fk9WREZjE2HN07i+LdLw4yUD
qKl3vE+Y3z/NYEF4Cln/M9Im+wZR4Ra5P9juTVIpk1nqSx+IIbTP8xzf5fA6aA1w
7ASgbXcHKYl9fgJ8kLydPh9e093cyMlyoKlcjVWyjx2nExSkZVCn+rO59mERCMvL
L8ZgpPUEgrDyW4KM+TlU9ZgvuwEzqlEcK63DooCiC9lPMlaRZ+qYhfLYS14o23eT
QjdnJl8L5/mnhzCJX5DnxsucjAsjgiAT7jE9KvxFqbl+tQxQaQ4cXgH8WEXk5dWw
47WAyhQDeMdv9Z5rYoTvrzgVUbl2TnN4WhgM0rl6tEBhqo7t7n1fig5FLfZ9IsHo
`protect end_protected