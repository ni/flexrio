`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 36704 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
DcaI24013a1ntsbbicG8f+s4NNjHEN/cyl3zfi5oeKGQS8SU4nH2jh1GHQsfrU+B
ByCr8swJWiTIyGxLjo4IZlyr046ZXMA/dDVN74eNNXX8J5CRNUTfQZVIqEw9KkOX
HZGIq7BR/5W8zn9+B383UIYlB4Gz6Plk9iut2bv8Dk5z1C3jvQMWy3v8PMwym2s6
iZs6AcQ4oSA+72DkA6sHJk+vi28N55TimjkP7lsP8MpTjcnAxKlC6EMniI9QWwrM
jSwWuJVSbikwseAZhrg4gvJcL2diK8m75k3mbIK4PZc+rH8t+9vowVcP653w9TjV
36WEtQ7J6At/MajsCxJ7d6rdl3hpcudZ3LwCZehDrbRaNiNQemDpmss/aVAAg3pb
kUGptI0YEGjoTMHPEQ5BrmZOKnQVaYwUfCQth/LKI3/ozxUkgCnpdq3ehn3IgLWH
/KbMrIqrQft4SdsIpcz1Jk5ouAj+anU16gf9m6ofp5xLZVHX4RKqJwCxKX0YDwS8
3evxlsLE+HlqY+xQ3FtV53hqwOixLa4N+WR8lDyWvs4sz2G0dQm5ggwzfTSEmiji
lGggCO6CqQ6GmPVOOcwA2Cskkvhb7LmnB0Qq7jKa50HHtP8JzwrsAJLoFUv2C3d1
EkhwR+pu5grFR135LDZpKZuGPf4QJPu3vFbOyI2z+NY+kIiM29XpCi+00G131Iik
VC8jve/dyMCAuRL0GLEXscIHucWAwlMhTm1SSlGPYAxxiJQE8+F5EslyOWyCRJ9C
tV8yNDAtrf7XJzBtIifqHo1gxhCmQxdRZJqMVMOAFyK2Z2fhTqMUW9lzJEx0OUYv
ISaoYFbo8WJNVWQwtjW+HX+IxYcjtYTOIqXaAdmGvjtQQNr7UyCuR9Tp5xc9PElg
xGeYLLkf7cZ+FyKSzTdqRSBProErRPNiigOCI8prC91UFlFYBxxe0vcqxYfLgiXw
f+dkFR4qZD7fsjBHO84A480mgcR+3NljLYmO30e98lnlBpAet4G78Yj7Q3udGzlH
Inrtsm7Sa+OIvXIHB5tkgRciaQpfY48el4ZahQfCGfBAbQSh/U+Mqx/paeg06MLQ
TSlHSCi7VzyKS/ifUt70XbJhH22+yGnPh+c9wx9tl5nbMrtGfGzxchcltNZn3OxS
BVY9ln0ro3OI1PK7vDtxQlEK3opjEepR7dLao1RHTNB1SSgUxRuzZ0AOc6s6gOwR
0cKm/iylcgojdzUNIxSmLffHHlVbNdjrVYv1tYh2zydpIhWP5ObE0NWgL+6obHG1
nvHLYPsbM6cuAnqUyJMTE7TtD3ZG1OkXJiVKf43Fy136BKQXz64VPstl+w68OvdD
LgVY+q0lq43JfDqNgJZ16VnYK9qNQwvT6KyOCImwk4hIrVmJ/zXKexdfAsdqWCFc
nKPEqr8FlWODKPbR7K0dSbdTYhjzkkw4H8XTtmBW8zfyWVPGdVHgQz5SkZY4i70f
O/4kp3Vzy5diG6QPe5NhyM7941HfDNhVd2+t1YjSWE8dGWtdCz/9nWi9ZoySIWJH
ywWp4654U6TGXSMes1yZAYA5Tj35FcVRXm2Apbm/rlHahng+dKQvtsviDqs3aOLY
qVQ5PGbNxRI2SGKaxcW156GAT8wgaoyQPaocypFRJH58TFfFaYiGQRD5b4xdxUX/
5BQCCJHIVmH/DVX1zXZcYdbsGYJAnhsAyAvMAR1rtuWnPrGdmXBymy90atxQDP8d
DVE5gO0ySJAobheWfLsaGymmNRVb0fZOJc7tSQ1mUq7ZcjPVUXgfRZxkEWyrt6bO
1ec3XQodnt/v+OfO07SnBZf78dnQ11Uz8SA9xaGSia7Whp3X1izv/HfjfwBnzMCB
+4+0DwH3KcHShJthOWdphE+bCP/BtIeDT4h/zf3du/ynWZ6cPAE/07ZAH5o8PYBw
jFvvWatzzY+r0ZEBVDP2KC9HMB/pZZBt4+VVXeXyPoGAd0pW8ELZ1PcavPsdt0t1
so9flkULGFg92rlED8v8SLoXNAqmzkz2FBEa18wdZOb6x0MFboy3hJieohlUq2nG
hR8oEcBeVjF5GK+NzZKWFe2UahgSEvlkt5+xTmWXJdC3GxK8bZ7jponUt/GcM+ZS
UmZzvleJRQl2lqkAjJVArEI09phIwBkAmm4m/4/pVe2GQ6aCFZte+MJATHxdQD6O
yiEmjbtI3xDtYBI7Arj15UVuA9NxHbRx/U9ojasryqErFtDHDq/6ITX6F4IZ9W2B
Kg6hcjHRCdooAnKoLxAuC+I5r4h4pxcC/0UXxdeBsIZpXge8zny7N8GdcBJ/rKAB
WnMWBt8eREFV2y9i25U6eXuOQc0qun+GIbl3AHMjU0SslsYsWce2G3+FDT8O0psK
mpF9SrPt/XVVMdkzwp4U69jPHU3SAMHXC+lFosOTgRj0A7jSKyqJ54VuwMCLgeY3
0whS/5dbfa8W5zHHpRInVyghIkBMuFFIRTILHbIRf8lsYdgBtfpJVmzQH8iqbWX7
7qAjNA6PRPVS2ZpFJoQz/8Mur10P/e3zgIsZ7Zfdl7KS0b/uZAVJoJ9G+igYTNW0
PG+1NxbbEuBVImdGS1XTLtMFv42BVmlXgPic7Fn2pXSHPtHmbCP7By7eJ1TVcmXM
bLhD2rYyc8J3+kqcSmJ81XYGDdhXL4Xj5J7UeB5tddODgpBWcJuE93KHNQF7k6Gf
vXS45gpCHiUnCkehipBZLIPv3zoze/bmokHi0CVX/DCcpbruQKdxHlbWzuA8cCs7
aQlur0Xcz9UahBkYHoKEJlzvPQTN8f0Dinv10CCE+VV+/KDhjTny7kkLoFSo8veu
AC/TdhFFJwOQa1iTBQl8GmmrWuBSeSpUo3YfJRTmRoYdR2XCUsA2gwbTfz+p++yN
5EkWF8RRwApvOYz201thIM1F4EfuxC/fHRkkLMbQLCOd7MeenUL770uAGbeODi9r
45N6mhe7Yhu1s1fXxm1Wwmefttv+Z4qfnjI2gIx27FDQHmwfHmyJNoCtUkrTWrNt
770Oz9V+GkQw0yUYxPgPj4JgNBAc1uwJPhK2lORzZed3UpTS5h1aWUQ71fLzfY/w
ZJLXAiWjdLhMTETGvCP8OV1WUOUbql+qf6TZxcN5hINQHlHB5JfzORMDW6wR5tTD
zun5ZqBYXhL1zmps58t7Re9l/s0GwmYnWfp5F/p43apqQFXJqfRtSyVv/pk2u9WE
OoJY5+/JZynVk96jd9rL5zR6378mhaq1jnn6gAdxBMglUdtoyfXhXNIIQVnkqIhU
CbYMpoRYu1tZ4eAAfwp4X/0zEsVI+WY0VpjQ8s0Pb3LRrD5ubYgBQvlY42pK40Rm
xI9UJTcdSC9++n6lOLbbqZC0aeAZPu+ZZdRroVie3PxAxG3q/UURqa7hGaOeyqDz
IC0HwHPLZ5SSdw63zxplkjvfwbfGV+nA8RUwbu01FuuLCZf9EoZaQ+CZdMQ4PGZZ
Vx6W6/rY4hYg9MkqtGSNDwoSF0fTnaUOwpG/g47/vx2qG6ZMEs+56iwnDcUVEd63
VS02ui7yzfudDzeY3FU9vwJuusvz4J8pDcda9kWT0nLvea/okI1VgrtGpwIZzvWB
dLtbrTsmCHfhJH3P4IFelilfbLu1Vx+7DE1FbA/t9dTbXtLP6TAz6gK2tapF2QhO
4ycKyOJ1L37G7oBZndFGdGtCAy7Hig5S4yoVWAt0VLCeARdHOGdIV9X/lcTN8aZz
6tn9fqEe0S2g+W/qTEkhmNzlzRiqTYXa2xfrKgx+07qAJGTpdKjYvPhd6j3/LkYV
MaN9IQ7HwnuZs03B1ikclimZxndFOzyDU3ilKj6se096fFzN4JyMCA4uMg2aUllt
pDoLEZTksNCvhbBgOCsPrKz8PW/VrwI87lwrPH93IXe/Ucugnui3qszf06ffYLUr
DXE2tUJsyZiRMmiC0S52BdaZ1mgbcfS+3xFbmamzDwd3HJr3/H62zmqONftdnxgL
9JF/nVseZTsz4c4JBIezfVZxAOEbr7ftWTULhQIbwosnCT2YbKz3aBtCwCjrIems
FbMPUOxcpHswNzzaReBQEygM+IHCmgesbvqdhcOklYk5u8EWhoukLatyPiy1PI0t
tOGV4VvhagCaOBsVQK1NTHJYnqBcr1O0xR8zomMDEu6ZdhZZE+2mLjf5Zd0SRK3a
32mdISEBc58gaWE07cgoLXsRx3xmuNzwDSr7PpX/wkmY1L0OM6myEJ42ycy2fgfb
e3g6XOvbbIBTFJD88ZXbuWhnmU2+tMDJU2X9JtDUtVgmYj77O+ywPiuICceSvlTp
pIGwUyVze3zDUtIyxwajgRxx/t5DcGrl2P6rq2FOyHmH+zzAGOLrYyC7pV1jve3h
CaSir6wA3SLmS1+VzEsHWIk1FyVNYQiHED8O2lAjd0rUQRSV2GWoYCf5NXp3NQ5S
IM4TyvOHcrQed7w9e7I1+a/6rvJXSi1xW6V1jQAOvRFea+QtIdAq4cq6nte7nSgc
LkyM8DtCtRkn6wC24Ti8/+Y5hSuTk+IBFZxS8nZFc+f/Y0KIt+/1RxfB53f49RZH
yAsHKH/ytUA3gNOsXgYEIJRPTTqZivIZShtGwAtP2QoqJv4XZZxsnIRdBxd/QOS6
MmasMx/tG7XM4Gh+/vAWK74JUUPZPOIKEX38/SoAHw3T3hqkBWyMSju/fCRC3NJy
CUq3TsbJga+bRG7Igsow2EfKI3UHyYF7leLaOWdZ6dUrqClFX6C4n8fpE+lpml1K
vd1hdcgQIiRJyfbGhsLvOkLDMMCFrkqxQ9Xmx7m88Yw862KrzSLB1ND+TwUbH9hq
WHZEtoDkxYBFf76484k2tZBJI0vxkMobbUlFgvgdHi70n+Qaf7y/Lzr04S3dFQ+Z
syRDg8Kt6iE+N3C1gWGYqBzFepl7RhpNX7NdNk+cydZKUT1RGnAAZtFWwOC+spzq
tPpZiAkiQsr4fC1Vm7ox15VRvtzd/38TTw9ROBq1jlsCwkPZrqPT33a3ugQ/tUDM
fO58cdjhAQLpxEWpnH/CFDphxM6Itb9YfauTlfHy+8CCrvEY1yD7PL+UPE+WQxWk
uffDGjFP11ZSGfFE/VPR4m9fURl0nEN8bk+GyMyxw3jP493q9ig8Z7I7zslZDuyp
+a/W8W6n42xLSxwdoRyIPojLCb1Lq3snikNNU3XGYcMR0MLA2WndRBwNC83F0v3C
mbqZXy6Eq+Jf2fRKY3N9gWzQSfcFa+fXx6brtf4OmD90grXAvpvlw+I5VGO0Klxa
Z9Zx4FpZep7rmio+6P9RYkiU4KYGAaDGMiQOJzQKPNztZFNtLIrWT8YTp1w9L20U
69E1x1OJFsT4t1UmAl5ktis5di0YsNuxgeLVZS8qDWShyF3DkbgO23ytKW842VLZ
ZmKPISJyOyhVp3X/oc/GKNgRhbQ5pCc8ltMZKGEBnKxRbohZWJ2/tSdUbfAkU6XF
SdLPw+R8KsV8Ppt3Z3VLxWER7/nOtwwK4zRWMpdepNSVIxc5yIyCSFV3G99NT+9K
gaAWkEuuDlYHFxi9VawSR1iL38fQNbR25iSjWMJVNSeZV9VJ7DEmjwCBbnjPetee
RGnpGwQT3oPIuEwqDMushslBdW3WLse2Uz/ULNbqJvWNcN/wiWmWDhOF3iJ4tENf
UmVfGOYg5sSIY5Rx1bL3z+vUSKrrvhBV2bRBb5/PulFTbeoGuGHXZypAAuu/xS7d
i3cAkIZVyQuwABuPS/dOYKMVVdtnvv3vUMJ9lkxHEZz6IS6n2n5t4H21ruEvaypP
YjsNNZCVrxv1s/W38ZFKHVt4jv5c/Kbqe6/kjNyswrBhBbqtIykrWsD6y+NOsqHJ
wfrMJZd8hhZ/F2CtMPl3+U0PasYf4nSeqy2quW9QKj9tF/4DKAmMTXYFXYB94l/Q
r2WoQWa9y9ZlKQjT0E30zTpcPK8o6S1Lzi4CwDdl+nbWMOEU22qus8dBLG5A5aNw
tPvc6brDpbLEChGEuEYssZ5Y69ufIy7n5DL+mGH6hLUA+LeAJTP/hGW6x1rDw1It
H/BeBfX10Ut/QGbGyrmAXr0+FPsJZO2o3U1IebH8owUoGFytPWpgwxFNSfDahmKq
DJEb2v1jl/7ZMiG74CXtSmhPgGEqOX0X90RzsfA3D3P63yd98CQcHlIoNKZIbmtl
E8Z3CPoZ02za67LgZscRCsqZExBDQBf/0q+WD9TL//d0vbKli8KYTuH1GN9/M7cB
aBC1ATVY1gOveVHzxi4KmqjUlj5BMn9NTP0ZI05CvRKhHFxAhxzWDIzQ/ip+MXqa
vW8WC28WcHIIAftcZ6h2sMveOU7qWoAQ4VlM0oYaftzbfN7NjXT0XWyo22A0UeN3
v8VH84AFswTxwLRrE59ZBVQdOFhNwmdhOayCKzJ4/QulKT+p3Y9cwk9xHO4G596P
2bd4NjZPz33Gsdi3FW4YB5wg1XF6m74VK1za00xRuZ2qN+5392DNfX9SQOLiA2Ce
zGeHyfzQ45nD4CO8Zi+i64x8Lf02/wsmxPQGmgDFwHP3Z/y0P5lrT5Y0e49HE84A
LXyfGs8buVSSajXs3F/jgbq1aXnAV5S1UDU9v4hLtUD2MuOaQQk7T/T5lTNFm4U6
TDs6XhV37Q87myA/nb8YtjyeYJn14gV3RBqhGCpdEyelF1t+sdsrvWOarHqYbdvM
4C5vwx3GxqRQdenRENF0RfAIjXFxMh9ConxNRkH46xkzPdagCNnzsHl68A0nhzSy
PxXZZDTK6/VBZYQUpo3vTIls55anZJoP9BSwGuud/A5+dzkO8sQHlklIKQqjMgiH
SKNp+Cn3gV6wmVU4UWHdLBPWuv/dAk58FtnF+U7ep5aMSQVTqTI+Ifpynk5JGbqw
orgrXsaOuCRLEb5ZKarhiXPb36ryKMvE01g4yxgPjppH0CfFoyVV38EHWVH04oLx
Gvr/O9UkroIP68kmR05vrTEvdLdHcq9iHnwuZIytWJvds0NR7sEEaseV6+XBLVtp
UhSWasTrpEQtKNmbnIdWCbN3KcAUIhxHLXvrWFdyHhRCcBMP9KR2FDJG9wRiZZ94
ihfao1wMaBIGVMCqQ4GkUf9K1sGwSS/gyNT3vLOqW7FvDbVguYFA2ty2t13IYCiB
Q9YcIYZ3NepXcj+HeaRkYvAuzmr/quDLIrnempSyKwNtyysJhEgJx7MUghxWqgrk
DjRrQUj8hiBNucWKDh8OcLq1QO2RFUIdPIvECf/1iZe/TcpEKJuye1uxt7Gn1kiE
5dZhv41sgf2nCXIOQ2Vs6DTW7bTBT26sICrAno10Dk9IlmO+4KfKYMrWYXXFJ4m+
7ah18RK8tuqCSZKTUpbOoeECQ9e7W91H4KL8mS8jXav+22guaZ7+ol7PNa1mjl3K
BzoVdfxsKcwP3XLTrYzpdWo/27N1o4elMX83Wv9j61hOrRNt1m1gEbhTAww7Dkp1
LCAZSKJfgzafD1juQIY0KG8EA3SxR1HxHBQZuvv8qlqiSRBv0PDFFFLeiIfTA569
9q8DjvSCm7Zf9dglA+NKo69CgDXxqlCVrLENL0xwduPZnhbqK/6bv+rRpDvTqgXu
ljKRPdL+m1zi4vXIuI1XdbFluc3e4+TYwk7C6e5q1mWyMeK9wjAlw+sN4w/1+X0V
/TLe7ntYV47JXeYNbflWPyMJNJPFOQxBKZWgdQKxcRY0nv9HoW5hYQzz0fekaFtF
de732SNl6jf0by1MdBFRRx0/R45o2RY5l+S6ZJ67tVIMgEmslwer2Agc/a9S6rra
5cyx26xPb2rb/XjjGJJQQV7SvZQ5uOigeXLAyryonM6W7y09z4ojQEkVYJoGPT3z
CPRZwQw4RLrKJ9lW9FnGLb9Lu9XHfTCJTy0ValasobVnCZILSW5xHbvw5MC/6IAb
5SiB4y6v8NUp432C8gRvnGNwWesPpvkBcBjN3xnO2OgrF+4+8z6ECnqKn9irt1T8
w+L+7DN7soOlYyvfWr6ynpPMoM8HBkpyeE3kjW+qu9MnNSIrtAGbR+R6ddSH60I2
GrVD1aAxhqTNNkf65ctr7q0RKy8cxD4d/FQhxK2A9M546/3m2/UToeB56ZASqjXL
ojCXxJski3x4FQQRL4HUUCHliV/kgtDDWlsytVP3snN1XCVNDMJ74ZsDUXuGFHRf
NFmDID/etZ3vI1ILPvps6ryVFnRqqKEDhFgc+GiC1mkvSwwKYfA36NZBcAOy5/ij
baRtXvmZaIlkxfgh8xjOE05WFaOnpm7foGE/V/2wPnf4dwGGDsQH8cL+ELgMA0o1
Z5sN8AwgVOoeDdnmq7Gi1f4p52R3wa0zLoE8HVfQtJiPV0f68IbfvVFPTkOVyJ/C
4Wby+dTMpueTAGHyW6nWqJVBPUz1Sm0qywOJFWJVUaMFWGB1MjR+4SMmWw0+cwWt
33OxOVZbuAy776vklafeD4szbvHfYCVIVEruPQmGKO5Ghbxh0QwjbGMsmz0HZuOf
jkdrC1AfIsUnZEw0QrejSeD1Rt2pogzWgVi3iU5p49Oa+z2hc0IaR1ExYS1BTQ73
05tenilhHy4DxQ2ihGf9ywiJQhYDTboQOZTBuJuiR6hFFpblJJo5TbZMP0sJR4wR
yHlicGzSFzK8LNd0o0XiE0mMWF/21mhEcH6e6tdVpU0CFKpndpEI3ISW7n69JeXv
8LieQAU+LNU5bP4fapuJiPNHEJxRhtWnIcjd82/jCTaV7bI2G6C+ZckAfrcNaWYe
VgCeeRh3wJQSDOBBVoY+t4LjkdpRsuAtIl1dGN2RYIqn4D7qf9xbo4QTt2eh5dH+
Brm0+57mIoO9XzfpADmeoCfv99R9kTBozF6MZLoRW6vlzGssem5wKOMzX7IU84x7
46WO6j+D7uHL8GJx24tBXUeg2AwHIcIwMMgEQNzQqsCkjbCEBJmmGz5v0I6Agb9S
oL9fT/ImuapwWLp3P939eMdql4msRvUPxQhqjQkgr47j4aS41ZyU040ZMsH08C/I
hi/iKV9D1miaTZZqWWD2/rQH2RpD1f9KyGCgPpffnPslYx6p38SXWeIJgmycjy/5
pCWjCoCcFe0L2uaAZ4JyxGDDjUg7zz9iJOV5P7FGSXWsZ+IRjtYpLQ37OQoKYifz
dgxjhF11hWB7zCaFC9+H1p1KcTA4t6vJdQ4QK32V/1lJCkZVuxKCCVDsnp2/Qp5Y
x6GSWKX1+XHhSoCOHmISA3bjC68dy7YIg+azXTH16Xa7NKAoBHJ8/vvelO8XNXES
c+KrnF5nVMruU/6+X6h3m7YKzkKPO/FA1Ja9W1tijSqDD3ZCOXx6fuoo1gdim4W6
xC03e/YWYmolbKWZu9/UbWPPeSSJf9EyqGw3+rCHyCZb7N+xDS6cROMPEPB+X3WE
cHcImow8EvkSrcXsBlEiIGwQ6tepJhPYJT+0WVHFFA4FoMrJvTZi1xyXYeGTYK5/
vsGen8XDCjWct19gi4/vBa9EaH9IzuIwSrwm9EfXnzKQ2dZTF563+037FIBfzMpV
SYWvy8jief3S967tei3ROZ5wqM6oDMqewVQmzs8pvyYvZVOL8fjrwoFmHvIxxcdr
Or5VSCNGIkHR8ioGINNleMUTZl81BmDh6QvQAkVEi8q2Yu1tibxXJ/rZwI2Bd59p
yf5Wj0eToq0Yq5wKikmv/a2rIEwIYg+3z1IzzZzB/hqXWjIFqT9b061U3uZkCJpW
ut84l04PYOmuU6C2lhEI3zrJk5ACHUMavb8bI5U3sHFswykvyykkdI3bt/nzPjLO
F016iSy7gHri1fJa1Gdlh2x3bJoRQsiKi+yWo8aTsGZur4rsQXNoWZtl2jWihiQY
qeRtCQPuWfj0th6qwNhRcxQ+GlJTXhjp/UJaK5e5nplzpbcftKjE42qfoBxG5e8f
i0OKDoYlBJuJAczQAUoUcyf6i7M9tOayfO/q7e9Ln3cMCXmafx11LptgQnP3kE93
G5bML0KoRw/hl+ph58fbJfba8dO5kGw1JK/2bl2TIIWPKDOpfH/4Wzw6eNKppfHQ
Lw1kdp+mPJsHLSvERkVqciYQJa+ahD8TRqDIGtwd36xZ0WliRKclVeaEQAcbA5xx
MSszIB/B91inn0g+OZIAfu/riBThiHaY/x3Ie3pLYxvAtZE3od0m5gpqgr0f1fQ/
iysQ1YQLSkHl+trp8czFtqJ451JqeOAASTGdqkbrgKsmA8mJHX8fVvb4jpLwsLg4
lD95WpoXC5y2kYRWPoHb/FolekUqxlEQ4ZCbnVeNRGzmkoT6yIwPJJ3vYqIWUI1t
k+ZVDx9qaaQeI4gVgfdtfGCNUaMQBYOjuF73bTJ2n4G86UdP/SiH5+5ix8w1x4oD
T02mZy/KDmaO3cjcbLo1cnBKCAld9j6GR54rkXxZUFwsznNJFqPwJNf503Hcz0Vy
Y9xIGSeTN2Ea/GIDso9qiG1LQaKYUycgOhxlbDLxncbmBm/QcRXfqDR+sN8bWXUq
2C4SJS90v1ry/yy1UYebr8lLtvy31DGgNLoNcoZfk8MIzEZ9Dap94urHh7ZspVV9
mfJkhYFg67mgsinc7VtyrMMZ44BUxE4r8yWlCHTor6sLhZ7H5JiSxYcsqb4VbGRT
6cuy2vWJkQuL4WlcSW7ESgfz3aox1rxAqPvFbX1rrLbV6NMSE/+/gmOFPzW57Lvb
tY9Jb4BpMWwuD+wJmNMbpMaWCywW8E+5n0Kc7E7nIQml+AOKfuskYQt9siCzZMmw
5r4VZKelNO4Gt9iOmfwOQhEoSxOUe2vnXCIUJBjIxPSWNa77znnUOD9oH52VXg1+
9wlTzpJEUZt6iFm2Up0ffnNBvbjss5jDVOTrvQoRrzDwtZ6qAiLO5WrZGlfx8BsU
Ka9CfDAGjoi+hhhOSImbc87UO+Lp3OHLfbRPjnMD5vDs8hYwWJvbz5VgjP/ZBA72
yt+1yOgLxAcmlSm1JobrBtQGO9/SJdW6mcHpyDf00eWxcmFD0S1BhujPQl/pMbs/
WBstlnl409wa1GV4aHZh42HfVOwaQYIrHiWW6jf/et29VJoxBJyVxUWBw2lZfzUI
2LQD3jN4AwwD1go6OLknoaVpb8lmK+ePrFRnQ8hEFxXcXghZ+E1d/SNb0FA9J/R1
y0Cl3e1tsNeCNDGuJKroeDfgPzxHaMRcP0+hBuUBwp5UbQIF+krWDH+3+ypFll9u
99xNu86B3sm/bzSm8q3SOL393JR4aT13aIgSPQ9EFS3rZsO+GYsNFL7FNJgOgrOJ
9M49APh7wgZr4jdthSZUFbKrrAr8uPYkoMbGHeEld9BBMENqWGcWodJDuxxnWsIY
BfEcQsVv0btkgj+SxGk4oOregYWp4jCYDfbJ8JTCL8gVnU7DGVnEozlaN8K5Mtov
RMzQNS46VxbZR5ynx4A9C54BeAuAm7uKzTDKpqwnJyTBB5xEj4NdF+2fr89N03HY
du4IJGeMTnwA65zeSbkfMHr2ujT3pfN0JqnIGmleDptqejzEVByb3mD9+jBkItw/
Jihp5l2EMUcb+lDpsOXjdqIunt/8Sf6mYHOabY/awPo7EdKw1dr7+xaTcshEh5iQ
392N7E2HXZExOibHQMzUZdFcxbxnh7BzJjJ+VcCE+3oQ7OdvuVbuIsFBQMaCbj91
KpLDdBFIH+y4duOUbCExO33RzXdPEyxLvr18R4bOVjVEfl0A7uCCllOBHMVtAThc
BXDInBo+EU3ofqaIJQ3+t9/57y389vg2IwZ5kSjeW0NsBRysCuYGI0z8l2R+p427
022x06kgXxiC5Qj+tDxLPVWV+Z+Aj0lT15DlFAPGjG2D3wwKosslYhKKGVajTda6
0DKQglR8Jl46LDn5FiWbejCGMwmnNSqMlGKg4wnuV8xq6UolbnhoW7+fv2h0sFu2
D+WhjHYIgQMeV8iJwKYZMW3qFyUxG3KgjlRUtQaBUdSeeGSA31rbnCgA6XnSeMUd
2xyyWEj3r3krgyUWOkeEiuIUo412WxOpl1ikjAG1z9YnHkIhEPnOpnJDO3sWwvzl
zVCbJ1MKpgEgB9ObbExM1Zcsr1GZ3AEj2CVFOlZxW/6/cC01an9ZFOCBKbgZAZOy
Um3f0QszWj1/LUDy8p4eMQ5NW/jdBZQD2DM9MHbHq7ufpoMnRYSY84UyLJAMJe6D
UVc3V9SSKmSaZbadeBBnfOBPLtIRcabxOE58NPEjPl9wr0ZdhRZQXPctWP9n5E06
VdUoYt4/MuzJqDuUU01lk1h+3DXJh6ESGdqmAbxs8Q7VeFiZVgcJSSNA+vKyFG5k
K5vE10mLcXY1VtXY1uPCuTPBc+hooW3tyyVNI90CnCngK0pnZnlBpLJFNTeh6OHu
54/MlXMqCtr2Nnbg6Ya+/4PDiQDhNmP0L1pusVe7GrxZ0yywOwlwo5pq46iSpF9r
kWklcr73o6llGkLt3rHHDc1QuugtOwzF4CKAv3Y6nIFbzo3B7lwAlV0xbhoJgYuB
YEu4k7peWw6iQpaayoBNa4sApt3PT2AEKdxp+zYEfzQFWwUYQUXj4YuIk/16G+bs
n9jMEMFvZQ3N8961ucQviagFCKfTZzbiVq5K4WT1W+PsP63/L0FXI2gmc8T5du85
ZNjEMH4s0+QPznA7XLMsIE/LNE4G4t2vLIabaa6MlK+O2NzsmSG3lUCtejPa6u5d
AlnTA8vJmVXlDvvAqrFw9I/f5mxR8YzS6kYo96MvqA3e/p6hFYkCpGLfaxGvKgtq
g/s5elmQg/6OdJpbK+zEMzTIoyoc397oit8tJIqByWZfYrYh2gm8rCTHu/igmAuK
z6pvwHa4iB4sXxz4O8FozvfmEWRrz1rOV9FlMWPECpmIO2x8ePWtKloU7D1pAuSX
uN9vYqeFerwcSAQukrWllB9zZ1hKNuCIFAoI/bVpb3VVh+dsRVw38k4iYT2RlX2g
he7MstwB1+OFxBB1n57CEJLoB0sUG4IFKR1sZL8kIXwBMAQxS0hx8XOGj9a6EFZW
dBsvKSmrnHeNmND2pTSrgM/juEhHMq2WIN2L0T0Snh3Y7DdEZT2JbPqovuTHOXo8
5qmpWj842L23FgDFxCNSrEpVxf+0u70fj9cV1OT628+eDj3mvh3sK/j6F/NlVevp
MfYbCisqltf1pUte4NUrqhXE1KRFvstKEsssF8I8HIpfO3p/AdSsz4+H2hoXhuLP
rL2Wlk15maXLl07bsolW0nlr8wDueUeVf+jicxZybJvhbVT+Vc8+Lij5U+GNhpzy
MA/xuPC8IC7yYIgk1eCoYnw+RsSY5fSWYnyj3W+udzIN3heqLA9tYIamoLxlHi0S
3u8KXSMcbkAUt1JiEqb7LapsoyzEhI1c52BFcXiU7aRGDJKckCK/3W6RqLJQJLGL
bj8Ykezg46PMUyEX2xZvg15o7lvrOZOOA5ct+3E0GpsJDpE7VN5lBMg+OfQvi3El
shqAnlNVas241Z5VsMPuOFW0P+j0JV8SgXwN8485mtDy6l0sI2uZ4+0UAapbCSpY
vB4Nb0eC8c0RCgvXhWBZhTuJs87pthZyJmQxkZCajM82HCexdEKa2FI/tl0+QcqH
a+Ud45XZcns6dKq2px5ogY0wMGSGT4WlapXbL5ZAc4qPIkI1/IM+DKUR7IY2et8g
scvxqtL37ypGH19OpZtvXnApvYY7AunFa02V53xskkkxzoCkGDpke08YMSYqmBcS
BJ/9sH9Uj8yJMxWMF5/SsBT7V1TCL+Dgq1aS7oFo+Lu/tT9fsGbPMmtGhg0YQW2A
foxNRnsr0EXWH9Pa73wQV16cJfcGcue2yQ3m1ZPVfyxdeTRLCKD/eeJBl4teWPHg
E2Kr4HWx7awMyYl160kzI3gQEpG6JZUQjJ30HEIoA2a81f2yVPCJ5M/RZ7BW1NwA
ZZxAvBWYYXy5E6VynWykOSuPHW0+rbrfANTzbt/4G+klF0R4lz8jClziE72+INz/
6m+iSLV3OhALtT++73ZU4dW0jbO0MzGqsGKmrNhS4ytkKJ1M453aumP3a0BMhmqe
9LIRBcmLmjerWdsAak+tQieDxNj8gGW1jCpOu7PkMPEeWG9L81eFROOjXjjIuKa+
GMvNzoemUTS/GIQMl49UNpSY3v/VWX9NdGoMRQsRU75Z+ykTloNUax93lo3pvaAt
mmq+g7MLbOYmITaiimP5aQAa/Bo3D0n9sCUOJYnEnRJ1wvxs+kPfIN3mbnK01bqd
PHMHakgLj9Dt21gbtZfFEFDuvrmcDwBZohVmXbSa1rjRknMZDgoMWVm3ISFjm89v
x6pyaoy+7w2oWr9E6E64PfUGkrJxruj1G+7AqMIW226/L4YihuWSnKuZN6anU3BY
F4wcweFjCx+YKOhbylH6eVNe0lHjVLjJeAQM+Ff2AZt/a3PfFta+vkz9ubhNfDyJ
vCTxmuyjswQ+C5TxeeCXZL20le3iqYwkDBu4LKMCLklPqRUDsNUwbJv6VaHp2FaC
zkI+oGq7Wk0ggi1zs/3H26uOUwh76ZhGv65iu/tyulA3ocnnrZgWL/5Rxpd2zeqT
COL1BBqZJ8vJW6v5i4oVq+KN2W74JZC8pWmZSKnZNJyxA0EUmDCjzBoz9wcf9Ev1
GsruBwKzcRGDqO7PBMg3kILiQY8MrOq2EkSurKVW9YdmTaGSkpLSLgIbvJM0nGlI
rsp7hskZBb/t2U0b++1JOmmkBDXAiJaeIpAQY2NdI2wCFLr3ZnD5Tr/SAoDyKpIn
G8FHUtiNOQDxQjPgnaKqq3wrdDL/UKlxhHdLutMWDeROGWfH7J+hPV2Bjt6DlRim
XngoSUP/N99l1t4OXsf51S0rHhg63Bqs6DT7tKqUpnxlzbJgDhBaRHB5QYC1Dl1F
SmOfoBm5mWfJTQOq5F5z1XUFMcOEtwCDWWDtAj0iHLeLaOtovGm/9f+lFyhKCtpw
lMblwQUHJ7SpAVfFeTx+vagXSVrKGcpgFbehE/fEinHbeEL6MPnDwNpq12Gd4QkG
cKtbcU5FvjBG7aAC1im2X8rjBtzwOHntwSV+cuHjGiXVPKbIMaj2KfXXO68uyOg/
1V0zsqLlZ3OumG2Lo1YoO2B3DJutAOWr4E11xM4rlFgUSgz4G9UtzR4PQ3vY4NHL
ku7asSd9hWM1HC9kjkAPx95TErduc6ViuADqWieWTjKwvLTxAfMAwaM1nP7VJmAo
W0me5lnvmNZouetk+aWIcV0OyXyhpgNNGJiP3Y36Q4jOS4DoN62536G1M79nxfUd
F55OVhGU7KES0Als7Mjv0XXfxwBZdsefTOnV5eqillUDQ9K88I4U7WNHbts29Wge
dkzkPdmHjmJS8c60ngpimjOybzDYRrDfshEJtor9IRLyAtbxm9lRNlKU5sDlbIJj
6iPDmStCO31FTkXoZRteOrT7rv6BwnymbOq/sVHMjd6+R5fa36RVk07Lmh3he3o4
uEnOGHzfJFnEmrtbY0z43K/mSotjvtlwo2m8da8zjlCqvqGnD7tl/n2ALhmKy/7S
Sch60KZf4LfiIYjDghLu5A7v/gBUyal2wcVuxICEo2d+FMdnempzE/EDWrRmiLs0
9fVw3PrLBdhETnoY2MlbyljS4gI23nKABJxZVy2DzJ8y7oBmsRg57o8heB5x1xlZ
aTGFprBejUs06eQQnn0gK4gVG+wDthYp7HYrKAEzvQpGTFLX9kIG1gsrmXYe3wM7
Znu3fK6eWtn9RMZM6OmrcSnk/UsauJK83qFepFWnE+3m62LTWydC0W4nrV2NoXvo
duyPolJ7l6uE897hT0jqmthfKeqb9noFZwOvWwTi6UYieQaWYc7+L0y3Uw01WcE9
u6dqExH3xOfktbKCVo/nVT/JahCCeeLrrZGRY05THKH9/eE40uExiz/VKI7WJiSM
I69cWCSVg0OkexYZayJkzRSccFEINNou3uZ1bAbfHJh2oq5wp20lwaLYvnbh1I7f
VP25Rc1F/lnV/z3KdjvUP32zYzYkPQVrtkR3uSk9IFmtf6YmgvDAjWo4MOFBRXH0
4xmFaAw9WXcuOCJRrI3xa7fqplyMwASI27iKXO3DIl0XDjrF/0gBUvEWGkaNqfRa
kbHte2eKYW4boPTh9qm8c/qpk+xlfP2mHACe/BVodVAphmJZDBuGJTE3e9Ndj0W4
8SFmUQOtU9PKtjAlUSQrO8WMJdMG+pjCqT8B/Q5Ehup+oGtYtiOHnf5BI8BYaIzg
fGjd1qEYspe+uuuggUSDmVpoUokVgNlxvGJX+1+UFhpuK4OMxRy1uD+d30uuegDE
JCo/H+PKTuFKG6KDxKcN5EQtFo6JrGauMwjDPPWBxm7Ya9lyx2cqbedjiLgGCqa7
bWvo1Ftf/BPHgIkydSEKykQTpmjMC6izkqsK5Xu6P9eM9LiKruhGYhb8+u877ycG
p2fcKa9WSxF9NrjHS4aBRrebIecXK+Y1O4DOiEMSk8CDw2qfd4MQK73E34xwhhq8
NZDXq/epB23ARgoSVnfbnOrSsA3xxo6jEEw7EewueJj5Hg9tvA4li3+lsT9MkaXt
SHfKAjl5OkPpgZ5tWjACfsy+XYnPfq8HXljUn01StFnBS0L/UqQ4jUdpaXPTAomj
sjErPtLZaHw9yVf3Q/YLFAJOw3XUyfK2raVxyxO9mWGFlNlVqRXV7RqcAZ6M88vK
U57tNiyhWGFREXIEv6CZ8mkDbltZ7pY0tKiK+sl7yqs1kpRpVe55+JhPoibzEFu6
nnTzeC7hfNNJYYcjtfUI5ng/K5oQOjsqd6I6FVq+RmaAZowbopb+hqZ0PHdHX+9A
EGVWLcxFeFnRRU8G1mGgQX5W70AglsYScSkWIzBT0K98bfzfbuZXPIW1J7TODIwj
1kguaPca9r48yLZHfAGjluCt6ODuA5l2Bp35rbYK6xbz5cMp/yrEb+ZTBc/0kwHm
B8XKFG0SiKWqdpr87ft4ljyhdMk8Jb2b6tZlydbpjvExha6LenHAmud7cnBpo1P3
DDwtEycNRUHpL3kzmJ4voo/hao5fiOFZKxQLV3DA95xbviQ5GvkOa/gqsAXh3INu
sasJQGrRtQ3dVV7TreZrRdYmjDG+IkA8X2JPgut5/VeWWyzBdxCvTxwU727FBe7v
j6/F5NK9BZYdC8EcjnIZ+6PrLxkYo0bwEC+pzFrjHOBvIfX4OMfsF3Rm/hAoX9qK
2EaJHypih0LUXgW71X910t0dZIk0Qv2xQ/jtmx0fKcJx6AGSEIvWeo7F+JjSALF4
CZ/WwN/+561p51w4joH4kw/91a8lX+Sf1iQ+7qOXp0uJyPTNwg9uri6o/T5HFc7A
Z2SOgK070lvAsk6qZEQ5+Ysop3/Bn/qk3b60xxHD1yCKUJTFn9kgPqNdopjN+w17
VymUGyF21Pvxq6K4qUPR4CVNCXUisOw56E/SvYnMg3PE0lC6z2zyQ19aBwPAJJqm
JAu2Jtr5/+4dyNB7j8ZE5CWPfDL6e9VrucCO3Oee3pasJILqnPYogNOjIBtYjGUt
8l9FZXn+Rv9z8QT6Z6GCdZE+UKjhLqG29o9Of4ABPCTw8ADkM8ULSWTbKEhnThxZ
fXtm0BWFOzILBcpnOknB3os1jTBXjXrT326Kyn8XhMGszhLBzhw4Rodz1leIO5u5
A3Vs1int4kevmEFyVx4W7JRapIRxcup8oTI8Kk6wTJzXN2PvvV+Qn3L+iRL+nBIG
KnSOUN2ePGjAwL+zj4W26iWCVm3DmhWgjffLqJTclBpleOehgjQCoMeJhMP4Snv/
A9dUdOUb7x+hf/7HkIzPKiCFgsg6qH52HdvT6VShynweOGEFJSTFrnnzCRo6YnkA
bDDdkr6UEETtdB7UnBx0mYJ+M7VZCEqQfjsnXf3IjpbcjDfDKeO7kmbUNJZ7hYrf
KnZ7A6+vohZ47RX7ZrbnhtFx6OZDVxPsXG22tT3ZSKgrfwYfj0G6vLo8Nc4BA5dP
92fC8sSjgvbCLKlUMNcszgtddwEMf8UCVEo9/4TZ6KPBc8DwsHLx/1UZsxL/nguJ
Cq77tlqxE/5KD71P3lse7fk5W3gtcj9YTX0LUCrezolstd8XsK2jsM9CKTvrEgEZ
Dwms6XRn3hw5vhOCgw8e6Et9EIJnoDhVv+cVQ7uGTXU5dP9o8RDwUIGigSwr65lW
WRIs3g7V3XgAeYeBsqu95bw/LDsZNkUHnq3WLLIDZHe11jYpnD2GdFnTxd7Y44c7
npeon/R+Q7xeV/gzjyBuBE5Pf6ULYqNjFQgqob6qcID9aENQD825UYKUSwXnYqn7
RZn1dwQPrLoe8sg/2WoZY+RUSIa+0rqS78jPCe+mUlGJy0dPZ3ONVvhsbOrYEgcn
70hvblcwVr3dvMAwPvzs0wUbq/OvCMCtgWEiaPicwlj0Huvyag18umODUVj7Fos5
SiQJrUKU7VP46xQTp6k7ZRys0cseNpoi9pkuJ1qF40AUu52topcjy6Trd5uvseGg
Av3ThD5pBZC8gElTWEkaOc1txtJQcI5+K3zOo7MBUtC1i2WYLQhXH/zb044ukhyZ
GDILvFxG/zF0EH0jI8kHeVDxKlom0X3XIRwmXxpe0z1MZsEC3SKH/waSma2kGJKX
wG+Q7C1DTYNaf7FZyKEAJ5s+IGSfXu13fQb/8FQpaGsk5acCUgCryX290cr3aAd2
GJOoB5zGTcNu128QxlxKinUeT9hznFhU1bxplv2e47Jzm21Qu3ZLaTt7vH1UA2Et
IC3umbdw6RYgqS8UxK3ldkfjFY/EAhEaaC7gdKPw+D8NntpFjgo91wLAs5oXbQew
hTjb658fIo3qpRvanYlfWHxXeFvNmK7uRAqpMu6V1sqdC5AA1FrSUVmlnXU958PX
nVd91Sk5ZzNaedkKCAKcxeiEYdUZhkVQBRHz5z6U2EyfXVIYazj4M+X0HsysYbl1
Xa9d4fmI4b5G3zaVG2/SFqgcTJ4+zx51FZQBXNHHSXW3hMW8ZbaiVFXjcwI6FyCZ
9zJTJTOGp0sJ9gMdVqOFQq9uurIHSjX3LlJFa2eEM/QDyPTlX7Vsin7vGMtQ+jSF
xL4l2yeqZ/Qqj/3hcr+Ig+95jlME+R3WDi3oKxM/SJZYHMsmaJ4Al+06PtppuFcf
XrmFFkRHSVSkoUP7rx7+O2laGqYorBj4mBFykdwiqeT2BkLSGEQBJbZsrj8aMNp9
eJ9VuEC9MhdzRcwko55uhGqEcXYUXBfFzekYm0A5D3yZv0DAIOeIixwdklAqCx4K
4X0SkMvSRwHW1xRR9xFzzgKc4PrMtimjxI4KTM8+wud3vy35EWNAZrHwWD8U0mxE
edMIPO71VHGXg3kmHgofscURKNVUSsgkanyUWyFqlEjmU4/izwAaOv9NvI+Li7tZ
DNc2CYp1aJLmD/EF3cOskg15YhBO8EMECng3lE0XdsMWGJgd2uXlns3thT1le2jd
Afmoz81XP8j1EjqvN+B+iOlm6H2V2TwrRKfgBUhtRNpgCpFkwYzmMAEyL0pC4Mvu
6XSDK77X+car2kb8T3I70S4gRMkf38OM4SPl2JtrY9mmWpCgyL8UmJ3fJTzCjoxx
uqUoRR3gOOsHSL320VH22D5XNODqh8e8da5czaRZ5wFiMvtpl6OhqvZT/5P6yRcT
+oxGeqPom5jVkjNmlM8mULaYG8GqrYUDcpyFrKM/F2S0T+eLajyYfROuXihMrmgi
nU/HmKIY8P/G10NI63uazjuFCYusNCW1OepEfXq1vDqLq28q3Zpo9LZj4hdI12yy
dgrxW4dUbRT4FjgL3hZdnMoFEzo7F1DWMpUp1yRJ4cCTvSFk9+0nB24ZMPqvXcpe
844nocoeO69+oHDyz6euwuTuVmFY5fk9z3z49gCKuLrCqeU7Ds/lwobVMcp7BcXn
cMo148umO7UivKRWuxCiYmV1WeuG7LvzZKw6/dCBNQLB6FIdTNGHIrglGQjz/gu+
qtfEjOjLsKU/s5aiFgvDr9vAIRLJvGHATJJXDsP2n1Lh//1O8FYNulCSTLrK6lTJ
PUxOPCO5FpPl9597Sofuy1CPFjbaSUmXwVlADDWTCdbL9GZUDSaakvdGOL2oU0zu
qZotRUlrQHx4giQjmP2P/zlm1eweOB1ql/wixVW45G/KPljYbrQjVAR0JQbTW+wo
KiZ1SKmA/x7t3LZOKZsbBdnxNbstpu/lGbEBxi1wd41zUmzHd80BpZExUPPQJlmH
2YDTtXk6nlZMue87idk2CiRgAuYYMqFIMF0JrzIxdlspfo3gftM68lfF6PhgCVFu
LrUbBjk259ZMBZ2ofN4Y0kQiZ+TbyRGc0WIW0r76+8YP6NFO4LUEwRcKZaPoZpRg
WapvdXBWd2cgA33fJo49ERmS14Kf1fsgZwLGgx9elUbA46hXgQOrWiz9hO+v8qGS
p+UWBVy2xFEQeA5nGwwpTU36h5Gt4xkSyvH9DQ7jm2lqLORV+FXkigwY+hW0VvJg
JzcSrbsGBxwNSmZoISg1+RkDs71qO+tMiRCv4uJHuUy+0p+uenfVCc8+Lq/EvJTW
/mmPD0TwXYHi8j8kfJ89sUIrGL6XQzcoOzNPC2eXUDSfmbBz27x5h453T5R84f6B
F8FGeKqUmY4ndQcjb4f3WCucC4YAHAXhQT/w0/omz+d+/OYkQ6rHaspR7Hg4L/ME
wFUqiYI2+nywLUTva0MiuPkAn1ttl8vnZLXPLx2IXYrr4hJviLIurB1pz6M7Klt7
lMOkADrEcWAHlwt4oQ2hlOS1iPGDgla3Ap6q3luAgpdeRZv07NF8Zp+G+jSKQpDO
qa6h+AdW3cGeWG+TgSO2yTY73tVILCcnKzJRJTjKLpP5IHfQwfDAT7ApjxiR+CJ/
5/BxNXMZSqn4zTQS5Jk11bzfs9pR/q61xV2FugL0s9TOweIRbJNQZTk+q7mAkznD
6dQv/WwSE3UFI0GwdSoU8mdIdNHSpxS2lbQiRBmXjPUYzvB1ooMgv6jMb4mi945f
71r4cwP7mh7AUhHeUEAhKleV8uXmDKKPj64EKjFXr2FnKy1IoaXSBsyeB1qYADQZ
5uz+k0o3McGpccibZThrOEnFbTKXOxsvV/laaSWWpn5EIPoAvMMWXhD+HaOtLHDx
lni/ex0KMbKcq6TNQJmGREgl+HSpQ+y8cykqr6LtNzbqJNJGDmixpnxzpJ9c8DR0
mEXLZtvnCS4JpWVf00Xj53YoQREy+1D3ChXutdd7gybyyQ8Sjv9WfoBTTZqcw7LL
lUIfX2KR341SQrN8PCqNvf+EvAzaJts5z419fN2n/YdMoCcNhGvV72qGFSYw/wB5
t6tqRXYVY+KVIuhcZ7YPLK0oWmBpdlt4l1i7QEtlTFhc7urgqNBPKo00UBffUzJv
AKUvWtwLV0iInsbNnwXMVLSrveXpAS4FjvLdXiJsm/NFLKYTqyvVidHmpCeOeH4W
4cvayNHsPjkIno2yFjsYGKCZfpaw5SEs5SR2aaEQm+X0WvfzF41UA9mWxiYURj4C
Qbj5GPDFWVu4Me8qTNjjq1ooG9J4fg9d487MPsu/Q4HJPdgcizOuk5fEJokk5L10
2OXxPFjCEk8J4G7qjyZgGpyjBjuP1kP03nVF7iVhY1AUN7XQtwhNj0Sxcg4zjpP4
gMg30kH5vR2ogWpLQoZOIXssIbN7WtMDZok6oo8wtkHLJpe6Pm0oKfjEMoPb9d+Q
tXVT3E/03HGCOkUo1zca3tRZRo798vfvd7zxQVBNYXKqF/4O9R/xpAw92A0OxeoN
rxPjucbZBrTr+oj7MD3mQBPMhi7wlKMe8YaC4MFbd3vz5D6dPES/SPhqQpWChRoh
HgVFp9ftPMdxDa9Efa/EUujPfg5feVJaKc6cBXnXN1iyHBBdUaLwjq/hcR9kFOcO
lExSQP30dkChYKYUt9Oyq1SKqZi+2RZC8kidp0K9OyK9cLPIzgS3oROiVbpmjpZz
/pxuUsi/2dcxMLcC+hSRTCplINcqCbKc8OAHdqpBEQQi+xUwn/Xev+gENngJM08i
RsM+ezuKcpoURpgk5sLwI6jQDncMYSU5ZaaPNUB3J8ECKWQkxvgQD+jboQRjwOd/
XnfJDDfhoaAQoNO6xOMJ/hIjp2vReS4yxpSBmS66wbY/I58Ve+xA5Tw2i3TuEN6g
lAae2+BNhMYR7vTEckh9IT2sVWo5JKwMU4Q6uDjbBRjRzr0YLbYhwNOiNK8TY3xr
OxNFyTVMriI1hEjTCRQT6w569cO2SlgQ12YkeoEfoVctHkzg2J6AnefFo3vGO6zC
L0d9DZnaDM3icT7PRp7Fifh0ho/8XEIxDuD2HSzm+15UnQpF+H9tY9s3pugkg8r6
ylk9aNeOHZB3gahAvhD/0RT1t5q4ZiLoV7XQX7LvnNvg2UJ8BiOwOerKEZfZCXJQ
YKZILFPnndRTKWi3n3Q6yKbkYNNPGhENhzei/ZMiElRhvbEEWYjOE+M182eI5AO5
7Sh+jyjsUscLCxp5WHvVdszWXxhpYhY+HkYavddOcbGG6ergHH+bGyUSxn7/p9JW
ExWmpFDN2RIGNLwqEdRJzoAFywRQXmnDOboB/W9IELfHMFnkgj1tWSVOfxpCSeIx
RHytdA4jdAJ8eNGcIccXxYo8sqs8q+R9MDQ+0sx3CD0D2aCLTno5wXpOjzcVkB1B
iHpnK8kKRoKMjdk36CRuBA/9Z0qRK21p1xiILjqCCTpwRmy3redLAPxHXUvmPklp
2V8KAtklKQH7EspetCZwtbGdwo7dEB3BlNCxSJQYM5qfbhH0CmTg7HGNnw6rDBs+
mBDS+t62y/S+gdBub1SrGI4oaTG61wb6XNlbomPqu4+HrWgk+8mgJWwmsY4BrE6j
wS2LnWJIbGAfeRqPGbYYFB5gxD/7DRtFbjsucW9Tu6Tn3iNOBH5MUML/btGtEvWE
Sw+0kxfdNxFqLnkD7BEUy6sqA56lyjdgxYTw3AJpQYod0h6yyAVdyFKGAGn1w/Bh
rglEIAonKtAN2mojaQLf3ZuxQxJ3BH4C2ooMdbNC//n7OlbcHE0t2dipBHDXRxUh
aEx/aheANZ1Zk70+rbHQZ/XGsHfeJviCY/Fxwbc8PqDb2sblgVzFu3q3gLZHnRJH
/t93YoWGnEknowM06NM7Z1iZofhmOFlb4/TE4gsjL01/nGo7IbCypPTZFLKCfMDb
6TsnK2yw9v+NuJPH0Im7O36y5ECp4GbgC1t5B2/zt7s2BFi1he2yBTUYQRxjgg3d
VaDMM+7eTbapNpgbKKVl4WsjmxhxlbDAfkR6XkA4FKTZY4WpiK5QtoowjfB6RyNu
Efna/7INQvkWcvxxHquh4EQ28KRcWeAw8OCPtEdIcpzaJ7Zq2Twd4VOdHGHmE00e
16RddYbFKtr2zIgtVIrAv4gFHy5H8cj/7jC0Pd0EzztMaQF3gyHbcIfN2SSkwHRm
/J/yymklqd20oSgAsEfT3jqyaBJC50CqP8UEbwX00eElcKw67l0r30B5aQAisPNv
G86OcY7ZXci3egaTtkaaqazUDLLy7EknCiy2ECLZV2+f0XWQQA2xU7WXWPE/R//P
cwggQ4jnkEnTEF+TKmpVWT61NsMrG9o09+gp3OTBrIm2DUd2ta5RyzgmMiLRS7oo
/CJyTh//KruTcWQ5ZsCdoNMg0ytUY9raxxRNR3rxtZET/oW6m+5W5cGHo19yidpb
MGHP40kTWE4BQuchsqFuPe00iFnOXaGPuuioYZMzcWy4xeC0VIgHEyYrF/5V1EjK
ZoUAKtOSKlJtavMOzcbbMovDvS+BT4tLCYCWioLlV3MN3y3WyZ0H0imXLQqJecjz
IIMFixF/EvDgH0DBz64HKmuTVEqeg6JXUhhB4Kk1Ytubq8MHvFAUz+rDRFdOucXI
4G9mkXghS/QsZmvbfqGdvGBm2/3hpm1PqjnOkNhhcWeCQ5PBC2xyQxbK0XFHBc6c
Ta+G20D3TZ5vEYRI7zk25AkOLMM6Gny67ROoE8/qgCiJIgM6rMXYfDx2lzRtJHYo
A9gdqmX9XjVH0F5PfWk1TQJE6Oo9OxRq2kWeNmc8BFkicLSOvhTb+YQvJw0LrmDS
XT60E1WM/As9sUzD8Y1fnKSMIfzDmk4OPt24QzV6c+16QhBY6qs5pXAoRYjfdFtQ
Vn7FakT1ZQPgRCIRk4C64hy/j9S7c8Zmtmh6x9zkNeE2yutoXlK6M+FvGcVn3mdl
wLfnwhdbafgVN3I6VbTpIShA0JY+uUMIIl1qAVTvCUJNOb4904SQV+X8HJEAOPRG
sLfgfARu6ykRTMpgc2RMj9wsPQ4kS2xKGhTSBBqMnburlAxrzecLrTBGSvr062Zr
VrU7OaXO/viEAV7rcWdXEBuCcQte7eNd3/0Hx1dRuo8xCDaN7F4mnn3YN9jxHQPQ
ybbVk34ZzyVlR30vWeXHtMp7HL5QA0XCd9CAwBuizo1BvC/Yxrvcm2e1GVNUFTXR
e/nAnBwp2HfcBANIoCVvsnJaQJtJmQ2nGj2/+2orKT3HEj4Dnpx25N9em6Pc6j/Z
sFkrTst95zfd0A1hAUJmUWA78D/1JM8WQvZEWI5k5xPaSnby5EmmMCmV3Opt/1pj
cViTkGKKOQJ54CNkG1hD2sSlAC5OWMGaPkF00QArrYimipUJgjS3cttoVRlh8dRy
7vn5Qf/EMHQvaluA0W9JLQ3H8w2BoayjSz0Dh2C6FIENNXqXbow2lq8daRbXuOfO
uuyfry2NYsqOlvJeG9wA8lOqnaCBsB3wlPZxdcvTZHX0TRS7Ezbw8SJWar0PzXeQ
/pcC2cRzBPW4KCFG0IPa+goO7GZZ6gOyUET4DFUVpT6Kb6ntnFKyP5tiAKTxU4pD
LhhFB2mv+ADz+Itat46qvzYQQZ4ZLw8D1/2pfCeY6TPUZqTQ6beuD44+H3AAmXXU
J8J/laTScdrZdOgemiin/ioMkJ0zJ+skj3eS9wOlmrEPw2vgwZQ7zM6ruHu1LD9Q
DAWdVsQ3d3lFijNGVitOQ0WN4Z3ZMQRFpV4nfmEwsILYbgxicDopA7imwFbO9P6x
HOXG030cEKfOJHg9wk277hybRTODUsp+LhiPI/DpO0G6gh9QlF/V0ijRGs42PC0Q
hcc4xgrM+B3vuVsAZDJS9IFxrs1oMgVZq1P9diJ3JSU4fJFmneJD+QfmhNMt9rXf
zMcxOib3KiOP+GfABDrQnrAJJ7GjkmAq7LjsagbXH4NPVGa0uLDnPVRzHl2MH5+V
3g9z05zLIOyonIcZqXVhY2kGn9fboFK7GG2KmcAyLpzcvBVCgKQe0PAuafd+I1Mc
7r9LKZMCgxt+35oIKoOZFYwu3WrXmW26N08rw+x6MKZXPryERbxroMZzl8cXIBcw
WMOXTiG0V/2kmO/BkVh4yFPp/vn6rVsW9AqCyqAXKuyeu6vy2c8Is15BtOPazbH/
6V+SMwME+njYy/Q5AYRkLaLUZgZ6l82tHvbD1rUiDa8mIWJUyBnT0W2EqpjnURgz
npno1U5oqy86PGlwYugtsfnX/nl3YyMFK3xFv2p9MQlLMZr6RuXa7zItkpFhlYzp
2MlVkmaJaB15JohFB9ci6nE9Vo4oLluC18bzlDeHNMhRcDwp1ae5N4VGzNUwpdIZ
9ZsDUztJ8I9SvOrzVXNjF2EpQgC95wq+FnJALgtyw+85ergp5zfLgLmjpUnMS36g
b1iH7MJ8i20k6Cx0s1NuIOdE6Av0kypRHQum8MYp4r1Mfx9KMgiks6/rK3QWTeyE
H0jy11Rc2TpkBAkxzL/IBxURbt2Tipi4HwuLFqDopaec7/a7dcl9covuvo7mGppd
pwkEiA3/78PJHFNZClc2MX/9mHCv945cUYB+l5rngV0XxToRXY0kH1YH+R41+LMQ
XrrV7bw7NOz/9N8RoImDJLUGgTwZYtTwSw5Grc9SgBb1zy3pShMqlqU1e776cgQ0
hBAXiib7XT3QyTwcZ/jhJNdee6R3rnj9iBmnlC6sjEl1WZhoSCrfnJFF0YNgLcPT
06MBqrfMlqEZTmnegr+lCWxs3rf16VgjIhvgxUUa34mfr2EGEvLt0f2turYpadEh
n8Tx6MUdlNJIEdC5voeOk0lJSgMWsUR4dDVPuElNdtMUwIPwVyM8XYDN+NpOmIP5
3iCGblFZ4w5W74ymd1UH/3AiJBAi0uAsfr1ZqjVy51VN3vkMMu/nij0IAfX4lfop
NbJGB7uDYEHTy/BXYRKw5T2Ahm/LurM6R7B8gqdvzknbib/m5N9VdOlXkaSXFoF6
yoQL+ZtwqNMXW3iy2CmCMM7dnUlCYZpZ6z87MDCKRP2kEUmGIfQnZs+zqRlt/WQF
gjFUd30dHZ/RVTkrYCcDGgelYaDFATapbG6dYIC2zVbs2arINSqyz4/rj0WSvloV
GUzwL5MYqNdCVxPCjxUse1OL9JitCSe5QiT170COwZyWHmMaR9AJcsXtHhrbkEDL
biTGV9vO6M/lQxqGUM6b9Wkc11Hq8swX9P/mY5lKSTPKdSKsWRmZSra+zougf2oy
3gktUSPZ5z6LJVFNNRebtB1eyXEdQGXCVxQc58ZrrRq61rtkQb/8ExUDeRhGH+Ao
tIExQy9BmM9D6GYxCTukIHk00fjVz9cZYSxRtbJf6qoE1FZrglrb5tbl4Zl7jezq
ht93mMka+jbctprDLtb2QSfkXOMs63F2LB8RvEHfLclf+VjN4L8EHoRLhn20izwP
o8jtrXDebqyMpbhXY1O6VF62iTmHiMWZF5qpw8FMaeMbciKPZqxN/p7kVrQXILch
unhf7jfBt6DcFpQbaPwA78zMVr2Tq3gIgGS1hzbGuNt1QAQ8skG4Q7Xx8wyldptJ
0k07FwWHAWH/zWEfPVGJEz9P0whClRG58GNFVJm1JKnRpUOHTbBnjIFz/6GHTT3A
cblqxd+szWZIoKVWE+pyKRuB+dWXVp8HzJT7diCaWYb8blMH2zoczq/g76qhrKkF
UAtRIqkioeJxoShyh8Uit3tE3hhzSfecgUU5Czr94IjSCzGD/sbQD2T2YPF0fdFh
7H6MtCfQchpjXNXo2hdlPWOpJzjt42H1wHRt+5aOeNmOHvRrF6I6V8AAYcoSjMui
/UGcALRHTh2jBm622w1MAAMDc8g8M/e6jZZmx6w2Ribmi2WvT9F3QhLajMlMXeR9
/xiORuTEkaULoMteNkGp2jmhlhHoBmU702alxqtUTcecfqO7KdOMHWMjeIhzNlLW
Nuaxyntq0drnqVXwW0qCkr3ZeojUfKi4VgnRnhPzoUJyVnNBt7kAXdEHGa+HWWqo
h+p4qXIjpecJ6c0CWdrVvsB39FIHgdiC1dt5QAYoJHYHpM8dzWsYWtX6Zyl2hGoB
c8DZXA8A8TaFM3UyRh+7OmyK3vfwjLEpTbofJFF33219oYwkZDme18OpSvGvDRxr
hdtVowyEAYRcNkA5BrDAfMOCdoVogQJYSh+GjclFuUIjUHdp0xQKlM3HvUiAz74j
wKC3c7cg6ouCqJVMrdGFa6BghLEOw6ZcE/fU1V/H+dZzarroUaCC4+oB3R9wZUbm
NaUyW4V4WyvgozWSsVS0RGfuUbIyoFfdIsg/bDESmVn6jbPUzk6pww0qQy9vsSd8
PYHvKirVmUv5EDeyVCIuBoufI4XExY4Fn2N5rYz5eKyJDAWY8QpTu5fcRETYmmVg
V5lpAlKVKKsW7t2uCt1gdQuxVYXvn4eVRNo2f0nX1kyk3wG8oYo1p2IEaWXScjq7
OjluRHKW78FT3FvJ1szcd1VKH1UjxHvzvgsy+3un82vI5I6/rqzqOCpnFfDgdl2l
PBlsBelToS2mhFV2hCzjBmvFrXLxrga1DS8mXqbZ+M9d7LaSUekaUl2yeF+jbKEv
r9slSMk5CpmiHtOxgP+93PPPakbiQ7WBq/GGrO8SiWUPBikqpRdzvRVgTA5JN3Ar
fwSHBN3LeGZAuuqIfXlIZCM6q4HCyEqbybf7ZXyzawZbJZMzNhbXoQqSmZxn8Ct/
lkCiTd4xXOKQY6gIXgt2GT6Q5ntBqMEk/a+XcWOeOnDfS0w9QSfdpOgeNCIb7UK2
k9/rDkVNA/8HkV+t4cJrvU30UOx/J7F4oAoUUPCK8V+ccMuGxdnHYES3OOaoMsv8
O1ZL5l9Mx6d/PL9eVH+/7BvWVS0LdjGUYY32aJXwDQtAl0SwNq3SYcTKvOTNKtg9
F8+fbSLsibttPZ2SMrXIUexcK5NQfVg+xzbZ8ZSsTk0eIVHr+8jY2b1zBODuVCLG
90gSs/PDIkxGLYz7qpnVS4V6lLciuKLEY4AzjkH4o2GZM3eU229bXK+mccPlpnp6
+1Kd+ZPlDOO4J9aHNokwyqMg3nPO5llI0PbMrUe9Ed3xXUzyYoNfln2F66fgtmsq
9rGmasdGUEPOEI5vMtdAeFGvmR8w1MoR2WqZqfIQW+kIfWHCT/gJPiezV9T0PUE6
6V1/4r823ukyoYLMFY9JuLUv094IOOZZ+eMzv5C7qqnHmXQZXRrT0isU+wGzr3ls
jRiPoO+3FGukurXYkq5v/MiLZ080RenhrBFBchZYF2Z4Q2RydUN20tfIT1f/J9Ro
dBYt9uf5/Au2yfQER+4wG6pArCWWoty3cUhvR03dINfWqap7XGUnvpcjXu2orl3D
ea5lxC2Tc2DeTKAkCahE+ugl7cykaQC9P6KSlGf0Shlr5yJqrUyZKvfrd/KumYrK
ndRZ1DiLYNx+09OvK4mvzf3Cgj4HGpQ8t9y/xwsrVWleiClMymt10kO1lEV+VkNq
KAdI7Z0oVjX4wFbrrsEBgApTvwvYaxjgWJq2erebjzxA+p7YTlAwPQwRo70gtV5S
y3+qvEqDKr9FiXWOaTA/4CId2J4X0ZGY2JKf35a30A7YInLCqiEofoFQE2MXaWQn
J9DiDkFIrcwbh17qWkTOxTiXv45CjXWov5RXZpyyRe2Y93eC9ruGKtgf1BeZU2s4
dOKNOEJsg2pGRIIM20b3/vMmhJch01yuY4qA0wdZHbxRz2QVpqIdu7EeaKkw1/JB
LvQkVC8o2huH/tBoG+ljnm6rbKh+IE53E4wWHp+GLnVxbDthZL2lBBxcbYzfp3ws
f4zIIbIMVy+Oumpv7c7g+uwS2Uck9jkrgIYiVcsD/+hgOyqaQr7rMgdyd9pKGVyR
J7kuz9ebUNOa07rIEWN9cxgYmG8XknnEGaP7PFccQ9MVj9huyIBA9MBYH3FGZbki
6v+tIZzMVWVlmq4UNJsZ+101pLrpRmcgjKnt86HrpH8Y2i1sl3GsLVfIGJj5wROa
oE/XXtsciy2bLoKQnf1TjcQERFvQ1Ex+4EGGqBbW8/nTkV2ZtM7HEjruU08/isCs
Q83adSFwXafuLKgFAUt1jtc0i2XjRMTCrYDbTNL8lMeVXoDpTLur+q1BUTB8Px6H
mqESiARqFVTAVML/GxDdWHI76A4s6teIuaFVJ3uObb55fzQttv6a4dGZVyxPekOz
EPO7iE9A0Lu+8IRKPkA65H/BmnhL+BfeTM1R2tbwx8bVOjM+KxWXyUGUO8G8tXUc
51sGXt34TuEEt/w3ViXNWdFjH+/n6i+8GgtwmSPA8/9YY5mO64D9n0ajWRf3qXMN
ztNk2GU0rK8D7IQ7XkkvFRgJGbn/hzPhdTsNTrjGcTc0YUxHq06AUhj6sLXKe8ub
mFh7lgC7lkpeh+QNX10Eee5zuWBYFeR8fXZtazpfmb85OVPwjCXOK3IVwC0LNRKI
9Hja9vkYEmXjcHzf5pFanzCFXTCLVh6hZYZH0F5mK2nLulGmvzbVL9L6LCkTW8Yp
gWbdgMyQ4EvpZevDbwXWkjntc+bywBywHYP3accUltWwHqzKTdcie7ilSuuofqDt
BWHTG3ed2SjNm4L8XvQb2dSF9RA/8wNtA/k96YFN2gtUu5VrTDNR4RFG+jkUHptZ
dFD6hxokhLK1qZcH+Z/ERwmuLzdNYR9B8gC7CBA97lAFD1sdTgswR2J2u2Cl4LSA
pBiZqTgiSLda4OOHDUpHCoXE1QB2j6ScLA9pxtL4VCLu6rzFhJQYEEnoQq5MVT6V
M7uvc4sMCdwEtakIJS8KAAzqe4PCtWeP05C+eiqVQKtL8NV7oe5kuwMljmPoUl85
f3RaXJhUI0hCfkA8WhAHPzZhNpKCRFQYVl0yPrTe3vh7mUgyY+Dsgctd05blr+1r
jf67b1578y2we69sjLg8R4AsneMaYR3qQRFlRcCVti1n9yXaJQsp87allU8kYm7U
pGIIWgY3FbPN7t2NusYf/j68nsXcOsQmoKT0bd/BcQuLcgqQbSuqHNQzdi665Hvo
k4cbqjhgwNS/LMS1VQTqzmb9FvfDQtEzSMe3qeZ1KqwfZF3s45psrup/b+RYxUF7
/vzaImz9RPl+ju3+Qy2mGZgl0qhy3o6oh4smlSsvFKx5sPAHPgP2hBaWQXj8YqRO
KbGpEggPZR34b8Jp4kacYkSN/q47omoeN6UPo/K/EUoOV13YWe3hY1z+spQa12NB
MB+xWMy8s1TS2X7s32ne2J/UKMA6H/opechSYw/fF8oU3QxlJ+UCFYFx8rWnuU1z
tC9CwChvimxd6d2VsWyjhbGG0XBP8x//yMJC23k2BcsEUkNVY6YSTnCJfknNQF4R
I/09AQrixcCb0gqNzSxQ5rY6k8Rjl2zjQ7ogKMMn0hnw3A/wqplTmEsOudFcZYZB
HkBi6oCpRihRUldgBPcmU1dP4KzxdwJMX1MTV3UNEUZEKqMke5FLpfbWKVdwd9a7
IZLgxlQzPsUtd4hxpUob1soIqpPGkABWgRiwqnuHdoF6xvxzU2WOZdPVqMHwUZDh
2mXPKgnF31UTBc9DP2qnNLm8kHSq3W1g9tNbdqlESS7cf7hp3mE8/euW2arJkO2h
0aCfAWg0cqFieIQjSUQ2G5pWEGddIdf6dHZWMnyvHMFijLDv3sqFtj2HCsY6Cz+c
TiKAKi28PcvuJPIXNtKiPQ/PE3OWv6lUGcH4eSgqwnldWjx4E85ltTWACBLa8Ia7
IRIEysfUjej8ZdQBJNI6jIRaDR3kcmztjqyNULB73vFCsCSMcGox3Bcxxb6INQw/
6crhJO1XICrcM8KKN0QEpmmVqZKrh3Ty2kubRlp6XQ6rwPumkKkTx9eZYLqKzODO
pVFkrHELAwz1Za++Lk5vKUaFFfzf3h85WlAXAgVu2MzE6uKlNzIcvuj15dWn1A9e
/V5kHdiNmMrAL+K3JFqgpYrE7Ekfi43tPTppab5P2vVZKaVtfADovQurneRGjMPu
jFoq5h9sXBj06uGM41+2xjSoYtJGGaR/umZ6U69jPNf3aFDlAQY6/jJBbuOJ5nH/
rHOno3lBOxo4YTbry0doVWw+wlNKkuSdwYyezgQlZ/4dY7vxc2obbLjYaEuIlRXB
FmbD9aDyz7tB9thoQZH5uhr07PO17IlPqUHOwpacYkPelzwIeL3FuzMyggj26C29
1YhpgXT6CbbIzPEDBHmjvFZAvxC3dlM/xfHLZA7qy1NDwhhqE7kwYqEuR25NeU7o
Eof0L/kiFj2zCDlH3NqXP9HmPPaYmc3BwKABpVVDqDajkPweiyqoywWa3gfe4ySA
TFKSOOsSwDUESxziVg3QnuiHOggema8bw2XbbusYiF8dsSeNCl7tnw+YRzmC0n1c
NthTLImVLKtZ4jqgMvzPil8VHmB5EI05sWE5HhXMmwNmpzmFxOfCjLEGaBxBITCv
gZJfgOTFjBxtl0Adb0emtfhhbiUkBAYXzbqVhgW2qu/+bjZr62XuhkAGDz9W1RXN
JoWYDMkHCcWmy2MWKBe7utmWP1v3mZz53SgyUGLc89wF10FB0nbvuS88vOCw+AWu
2UFaUMtRhpLPF/82ixh5dxAlN8WqdWUeWLZytrrtwZkNoxMUvC5atQpz5N8Cexdu
WtwacTAVMBwQC15h7PkQyJYD/KlQLzt0VzBurkMg4xOvS6HlnJbkmdwomfm7VrfO
eLlXxhdfe2rqoM8ZwWZA7WJKAIgnAcZNTOxHUc4MKTUuRJH3zK3CTWCgSGTXS4Lc
UqjodC996okv6170DbTy+wLu3OWu1qYvUeJaaR+uUk73p8ygn2d5p4wP8lwGZUew
nw6khFuIzgoRyXklI02uaH/g2B2p0t5ggawDKo5/t4+9mRwpgnWXdDU11GwB7vNN
mFIXJEAwfA3A1D6/1gkaaS3MT8UWbizhiilo/x/qSiEBX/CDBwnFkaCmsK52YDrv
wCbhpKwGi10BAOA3r9jchaFICscBFdOcYWf+8abDEchAevS8AKYh4Mjij3Vi2X4c
J8C6wogaSnSBpaCEkvV8aH2uAp6pWtDLLH63D0wEfCN1Ni6zxQOxy/A7HybV8drC
KX3p21wObP19NM+ztRO9RqCIAojx1YA/xl8cVCS1LvZbP76QRSV3IS5dSCjByCBs
tpX7/0rXCI9YmkYFokYqaaZHnFNKBYEaFIbrwZLxZWXBdzeKNwcNpi/tMavxxlD2
WRvhFrySdYnfnVl+jTbESWbHsL0ckZqy7UsWDi5jPTyOVf6TH5sbIPMmPgHOyCGm
KeR7kHnB1BgrQ+sE46NxsMCH79EewI4nT9OM9CsCpWAIEOdNBSAMCpi5lfNlCyYc
ESXyV4PPRuca0xK9kyEN+rO0QlO/9tbbS3Jw16zG5Y9M5AqVV0IGZ2cpecnq52bD
moT/sQ/cUhICTNfjCjX+4Dttsxe3TmZ/yB/a45c1tdRzg8njVibELa7hIxyaLied
M68JksYcV5PgP9qVVL6Oaop6fn3oqhfO8KoczFKhFox5NC8Y1amrQ4yvjNDE1H0S
8pBuRmvPpE37TyB5VHjeFXy3idKlKglo21G6rVPFHPliK/4Qlv7kfnRXVNEzCD3M
cj98aVWsHlljQ+Me10/t4NrpX79TqrlsQ2X7yNFtqQM4mjQxv/H6noFriqD39MOq
C8x/J0xb+srU2bGD9sT0+xaRidkzWML9H/bNTA/ryBxtwXz1QkysMTNdJur6Nfus
wfUAlfOATSGYalAyrhQxhs+uuvEAPuAYkIX6wyIJqpQyYpLEL0gAtcNLqqoJPy+O
xKu3JHHBGMIrcw0hz1FG3a0sICKVGu9wD/lF/C5W0F/dbl9MobxDWEoNAZgpSxt/
y488vD3fubBAcX75M/g+j1NTnKOcuW908pqMPo5XYriIoJ1grdH5IUzHkfoazvhi
iNKAzv9enkn4up1ud2SiOHg/WePlFpgY65AL8rILY2ZHypCQ/iRqZa3LarRKBogN
OfQRMhYvHlTbElRw6inlZ4VflrWOrEyx/Vt5K8+9ztwhjhTyMounQnLv/3gPm1Wi
p/fLHdHul5j7bdsVZeEdKBd0sdgEEaDon4T2oIqgt2fUuwAsuJkQHirNGFyg3RC5
Tnt6p1r7XMDS05z4LtbJN614vrIQJRdTgWoFodRFiCYO1DHnTEfGPBwvTZ77rqrp
1PIEQWNrC+sYtiXnzPGu8U0CUpis+H6KOr9momeDQfhrBHS91kPsqOYbs8PdY8t6
di+lo8fOGAti1YCKbhn/Gcd6GQPcchf0qA2kAsmOX2TU++bwf+F8RtSk6sh7s7h8
KSUoOqovNE9FBIxNTuaD5sgoKNcv+Wu+hszT5VkzLiVUbhAckO479BQGM6uguibt
wtYjkvP59fAIHbxjYpm8tU50a+Q7EUo4XhoeTJrGYVkwNDCNv+tyA1rrmwjXQHWl
jjqqDDwYqGUq40wLKLJtPiEwURv1Hi3kzDoe0AJlZWm4OIhmDohrujkgRuaPqnkE
AjvgISu8IPfXhmqZRrSvoNjI/YluSAPWo6wgVUmuQBDlYKAer11njaCtwNMdHzmH
0TTUSHM1uQJ5fI0wa/H61oj8GZ+OtjzgO4IVZCflcoMx1EMrvjH90fAh2goSizjL
H+d50/LVVimbWc3LkcCTQ5k4KuwW/7L+7M0wInXG/7IX3Q1rbqHDaq4pr70WrX1y
/xJn3Br4MiXWdqzw98AoO1QCAxHZP9UCLIU6AFWCRhwZ+RZsJxuNDY59MU/lRER+
6clhknVp02coqvNBkGt854WIYigZusBl+4pRzNjbyIHdmZBpOZDK2646x3c3NTmu
ooKPhh/L+NEDk+kECBYjxiu71dmOzT/GsmSr2S0BondOUQdbGYOjxvLeqHOo46h9
rTBzeXFFs4RNSyMIBM0ZF6BxxpGa2N4eyCsBsMbhcLUHrYjjKWdz1RUI+XQflqzm
bOdUnlPnBYzKmEndm3rmFOKeyVnpsqHuYPn6mlMwntFGu7Lmr9RcMDQfPbeLDTF9
IbTADVR/Hs3Pl/dQ3A6e9Vk2BNC5Tl/JzGTzTuGwjOIuUngz93j0gSgGEwQsO5qi
rjlByquZegvBznxSoSFHStvUf3R2eilE7jK5ogopmRKiO0lzJc0llC8ddc95hULC
uau7KnY8h0w5eE8u5Y87VNle/3WUBNMgAkoPgCnuOL6RF8ph2IcSarY4ZgO3e1s2
XryH9CbDsIwI1O5p8M51XzaNctsXLn+hu8s27ZdRIKmplpqbL7McBFoPAZ33tLku
t6skHcq7DwoK0YNu641507kLb8HS4k6wGBQsyjrnLpp2zBATK5ss/tyxxgbh51L5
no5TmG+1WxEZS5X3JGJxaRqYVLatssVFv5wRY+qb9rlFEMdhrBkpDT9roUhJFNqJ
gxVHfG6VZXnhfIjiRRZDrLP+gwNymCDJXLv+Qyk0GoW8z6U41cOki3tTsxFMWWkT
RlxwoNfGlqW7z1Ltpr+5rU2Rvly7seVAjt1MWjT/9C+epBjJM2OnOye/7SAtVmkJ
HS6FWrV1dtylau+nSsWoBwjcLI5Sv1ZPHX+MgdG9IH93Xf7LzSmd90wWUubXKKs+
hyx4xKnzMjBYJHO1mXxwLylbLyJCqThxXhJ0pEx4FrpI1AOLrwqyXu1N64mAz1jR
UY8vodtTJNMxY2+58jAUVMbDtH49+NMxwC312mAhQvELbjT6mRhQ2mSJ+tGFQA1D
MWboDz1qe0SGxDm4HHRl8R9fijcLBoVzc2++TmWSFUuwqhcVd/+fP73wKyYLTaj5
anpsqNoxJJFe/gPX+JQY61wfT2dGR/hyCajgu/q2RrltOzxg7OaefQW4eAQnZ5hu
b9JqdGfE6h58rnEkcfpXAm2/NCNIbTB57UG9bjDkiL3gxjuu/l/yxtSJXehgXtrc
S4tJVRFfPnonSoEvDWzsk9lMkues3sCd48VHR+xnxO/G/qbbO+O1FQEWrJJIFYJ1
y9Co4yJb+s/rHCFWlbA3SG2ip5ST9ErGS2P3kXeK6Ap9yai3e185X2C5K9rs2e2V
JVDu7sZCLALRavqXbG4YfMSw7BgWS4WFfnVJnQvjt6AECXpwxjvRQamcWFtTMLQb
YXxTOpp/WPRT4fn2i9kNP7lwvIRdJZPxhoqeasULyBrwWva3EHWCxLObu3WEOK4T
AQkxoftE7tQ4YmFs56CSkGgS27Fv5pnp/7Ihdcqj8DZBH0l2N6svmXbNMlmbxq8O
1vmu7pvkc6M6ekdPTcPXNdxkQLnjgi+l4zS3sllXiCY+UE0oMtipo09Ht7wZq26z
pi5ukZ+ON37PTU09dvpYhpzgx0RZ6Rem56b5A5iPd2HCxWhbZkTayWhoJMTZ0/IF
05a4Cpwjtk2Kyh8ofZYb8Xh5zGf8fldHlIRqTz/Wm0kXHOgz6FD+PMI4ykw4W+Jh
gIaBwG2gC5JtkVBA/KQd6SutskvCwOV1N++d2Dzy3LwuJ94YU2axPFxnZ2y5Sjy2
/CT21ZrJ8bQmemO0wekPKTdpnxUrRHKjvVb/bkr+v9nYpge6yLPmJ6o2ttoJmGt4
wWoLz4626tsgs3MzcFg79211BeVoeRTebWNXlm0jDztcNBDOULdd9AaMsVunzXne
/KgxEB5P1yPXsuhDeSv9UhrIcnd8cynN44zFpgHZA8G0QD4EMJJgC276F0tx5svp
SDuHcDWbrwJ2NZytxl4E5k2VAIpPY3UzD+Nq8SuXzGAIaknQpo6Zn48emxoye9u4
jynAq0HXUarw0GOMHrRq7UrQOVZRCwss74QkSAvm9NyUuYA8Rg7eyjLRQ19IU5Ys
aZEt1M8VtOdFWs7pInwtnhkT7c/fqRAnMAm9KSuMm1T4Zy182y6yp87G7mzGwzxw
8n1ryo39tHpP4IawP+UsA5I6P7fcmgyDC78ceVZ31+23lOX4ofmnefwcJFR0QVZU
p/OYpKKxeWe4X5oDCt7/T7njU4KqazRCt4uAcWbkVP8ZWRcs1wiiJBwqv6lgOhIh
vpZvkVDKGA6O1JCmHwi9SLEWmitrTzVqS/ZFVZNPtr7Y886dupe0I/m0UC/IP4Ij
918K1Pgw1IcLdALB55zilB2/cfQoap6Itp3EJktjCe2tiDKHiefFC7on8KsrMojM
7c5CNYdtZj4WhWTvBoC9Smhrt3BvkiNUU57dJCPeohopGqdwokg/LUbtQQiZcbVG
glFNAwQDQoQjliEZcgmWdoOM2d0h6yQs0uHCVg+vAr6IAV4Dw9D2Sh9huoraNWjr
fY/dFlp8YklPTMxzLAUp+CwtaiaQFMWpncwvpg37B4nas9EjR0CJR33nI1b7YnVJ
opGpoArf1Gd8JJwKyV1Ve43xr3Fumwm6eXNr/8gtG4ZWLserdfVfjHS6rGKsKrdG
f0adkoOit7xzne3hMLq6WXGMw/qdnysdmSCMR47vw3/oY5/ayQpP7ht1KwiulYCj
0fVMiN4s4e46jRo9UU50pqe2moitldq2RKeET9wPavCvpigjYJ9pxJqFAWNkwPc+
K1Szcga5YrIQd0dXIHDEpmx0fD1AWLaC10kremda9IiTTNdxjUiA+b+0e0Bn+A0+
tbDz/X9jiG4azB++h6MA6dvazsPZtNfWHqTrJWj5lQrXkNve+WVpVhQCVRMp1oul
cjXql7rOQga7EMhOMaL1yQXQpIE5Z25H145Foc44rJWUYgefim6kPB700769TbDg
Cqqk05sNMWvdNC2dgbJm4BAtqhBv8uQbJcgah2TJHtLxVE4T5G0f6iRk+t/2YwHG
A7JWHEWi3+yf0BaQqlF/zgvB9rdZAwIsJVxb4CrIhSP8aVPXSW4zhDMlkLL4+P8T
JHg8Ixww6hUZauM+86O3SH5GRZQYfsOddQq5f1gpAuKmDdx44ydmSHIQ0B9c16Ds
wz4bdoBAH5jh+5dBV8wonk6bR0qeU4xuOzesH6bJLAFJ3/1z0ReBPsPNGl3zG+EE
iNd+GtRQzlalSFtESWviCBEW8iT+otieKTIzHu/KRoi0xZQL4Wgeu+4x1jacfFuE
cSsRMpf6sGck88N8z6qL0p/sHO4U8TYeqCKs+KxHUZzT+QEWCMm4G1nYDBwFKo7O
yoOEJXSS4CWIuRSVnCB85cPm2p3NgjB36WHehGdgHCAAYVVgcmVbZ1nVTql8cx3D
BDJUxww3+8jtRKySiYeblNPSKNGgvLJ7LvfduQ3IiflHslfzcyztoc0mxhVXTRYB
1EB39J/vIbAn4Bxs8tqF+Jt7kvBxoXunv3p0UyzanNvV6y5UEUavus5XPtttuJCq
h8mPlmwmUbwdZJu5OvbYsvXR26q8EqegrVccbdTb7jHBIJcLZXUIMfYvAc829+I/
yD4DwTWH0Ewdjt50To1oegetmAkOncDmatIW80LQXQyzhulDa3G8kkxvQr+mQtO9
ZnNwcFYzRdeWPH+Hxap4Lg1xhTrm39ptTuHH3wjHMX6OxrtpY/IBF63KeOyC6GsC
zRbaz6RYUuI3PoFDaZHZFUTK189iUpePJujDGAOCBIJ+F49/t28PW14Rgk8hRqXv
k2zcPuHAiin/5DzHNxLJfBcgXh6NR8kB3fg2vncbEXK5jhIGWdyuoDtbNB/ZrCNv
SiLkjsmsqvEKBcMMocl+YMMVQqGcgfaIJaJrnmGWYsoaa5UWt7hbBaQ0piIu0b5O
dGr2JVn9s02iDRRMnk4fZ0HS9FhhZX31ruCwHNYXJaz4LbmSJ9MbEpBRA/sqX/7c
IIorCmZcTCLlfnI/NRU36JztSgORg6cV8z0pExnBwIT1uP6E/BbhDwoWOABBxGXi
3lPSUPCOO6IVsu7bdwWhyr2Rrvpdo47YZzwON/IuyFh+4brAxmeK0moc6ZnteHG/
IbosZso0trgRpzWc8U4NYGDF7yKbgyMoy/9eTibmP+XZwB0gWH184FKfo0xLKR4Q
r/vivyROOgVIzixqTMDu+F2KaAfXVjjKuMTYGLZrwDIE5xyHODD+r5BlGY+PURAv
tfzzzb8IVO5BELv8WG07yim9+jOCH8e7CyqKZO4enGsiGiHSDipw4viDtJkCLMSN
LDaizwJF8JqBTIrVwaLtXDS/PDLMUS/W5EFpoJG6tLExr1UHQMbidPwNvvv9/PJY
sjaCFUG3pMCMBKraDL/7mV6syIikWJBcOWn0zIBYmOuLYzMUUz6XvFGLmRt8Iqag
6ICZC3rHpfxBymu7oNCo9zJVHIpnln+QZpXTQcqJA9u1z85rnb/tStLxZ8qpYBrA
3OnkFBJvd5FTSaRJ/8ch/VzIBP2pbX62W3TQS9VLoOKNd627DtUUH6BoS0Xg/aB9
FJMFqrF0UePuc3F911NtVcYua2LNOw2iLGfxsKqKCN8UrOy2idQ70olDAqGvUvEU
/FoJAiZU+p6ucZB0Wl8vEbY1zB5120y3Uxf1BCK4jdYB3fQbS8aaFvwPFIh+EJzM
spmNrke2nyNCaDwYSxgdyo+Z+SQwgtTv6WWf+AD2zuGFcjbOSwQ/Akq5uKerc7aL
uPn0J6MW6u7K4kYvafyrLiugQEh4ha9WbAe/sj5fwGxZYbleOvBXU6HHVXj+6SRy
Z/wjr2H1fSOwk6fbukFWmONKsuR/5Ex3G0fqAnTq8L7AAZnPzCyhhO+N/k8WN6jh
0AhzA6E+L36ezD7Fbzcu30k2xcWC6F4cujgYly/IJypiavu0OtRDFqcuYvMZkB22
/HqWPHK/YeRgaliiIjr7AlzwybbZVnO+gOa57KA50s+UpYAyh/8xnEE/eVytIBqI
tEp7UvQYcu5Hlk9kXEIVk02Ve72cVCRUxGREKcHjoykD5/lCM9NvHTbB1caHP33X
1wl6k8EmQpWZLH3gfM557Un0WIiPen14hOQje7Zm93jiBxOC9nN/R9ujHYHObKrV
mIgq+XzqMrwbWmS+jE1ydQ7CtT5nnR7TKXN2/wFkphJpoOe+p1f2T5dST2epSHqe
WxYBbM9XJRj9tOaWqH7CauWW8TxJyC3K5jPrJb78AQ8mZZgXBNOYEZRydtdxqg8W
VmA/HV83edWLEHTjJQb3WjtSNxEPud3Vwj3/t4R+gRNOcqv+1Vi77UtPXwxd3hf9
s4v54IDsx4gM6HdbwnUBK4dsGX+e975XAefcFdnZmTPNP+ypPw8gnFg1bK9gmW61
GmkWGZAXX/t7Q0uUFN62F1JPjGf3N4hNBuNWnFlTmndpTOPkm1GX35U6PqUSHLUw
KupTQK1JmGeeSmci5qloU1fReZ/9JKlV2zArpg2zGPKrCS/fBqxi3jU0S3oS0fjl
6uuD3KCkVcLnCWJySzk1CDN8EcyBFxIP37krWHNLc/m1Vh/D3cYvg83mQDuI8jtG
b1zqFnlAAwcdO3HVFdB8cDtBqmpeXiZA6+VyFjvPMbLb90C9mejOg+LT3mj4JfRK
EZf3q2XB6k2vamqYh5SMQO222Ctp1llPTl9GGgvSZB1VLGI8q21I8Ha/ec8wda0R
EqAEY8Vhom35egeyFnGxklubr5tn2ssE74gC84m7cOUNHDOURsnMU30crwGrNnUS
IuC7f6S4ji6OvCp3qsormofHbTrxEbmq8r/W7dcb7829/6MFrIOJpr8ufox+QWuL
3B4yhx+rvNoUSde26LgIU6DAMO3B41fZ2yKhw87qFcg5ARdrmPsgXHPNpRE/YDtI
I7beafAoKAE3/RAvduGugZiKnGFwpBUCCp4SftYgZP3BMubi7u1oLYeVYTkKXxz9
XqWdDXzFGuyvPr7DJOHBK5swX6lDCC1MoE2L8gzsyleqCCo/lsAHCBTWFrNWnifq
1uxo7WQf/Du1nbhijWtMK3oV4EKqw198RnlzZUzxpfdCMqljUGFQtQNfBNKJoLC0
eft7sQP+ur3Vcpu740ZS/Km3CuEVTJ2NabgUK6hRL70Z06k2ha0qJCMdSAx24h+H
ojplXkvm/doIin3yqsQUOJJMsiY9cyXhfiJ+sKnolCZB25tm6x+4C7QxijYrDrcS
QaYPCeABp1q2QsyFeVp3rLjC5nSCfsirGLVEwOc4xqluj7bRNtVNaDcsZ6S/tlTR
RWJqsn36+pcVobwUCt9UCTwzqybxBkF2111HpXIbnHrNuVC5ar3B0yf4XK4q09Ug
XHRUfOD87t9Fj98sUpCjpPDMTPuh2XvDdxwTl23kqJ0bbrq3dG/F22q9pb8XV6Sp
9XAhNVYDDzO7xV1xVA2KWimaS+r2INrH6JQbnrc63fwKvEnnC4y85tzEMsqnnIAo
v7TfgI3qS5NfO5KDd7RquZK3rbVMwDcJRaYCwy091N5Hb8CFZaPsSOHoUTS3Daas
GzJHYQ+wYaIEZEAQ6HSGLpGYFERJ1dY1LPGQjgd+J0+TaHDILdxPxShMQ6o0B0Oa
HucykISLcY7gwRVXpelwY9oxe4w5qKQDSLcWnjF7+3CS0LuhNYjVw1iBdqIYt74s
DRE0UnAHinQJuELwYd657lvVpyNeyOAQqm6gZSk24qN/2qdJUaketF4NamDQLKK5
nCBR46fUPLdgru7tbxKMW23QIHIslFnGzWUcsrDX/M2XC4OMaZSwkYS24FFoqWpQ
zc1NrHC9a4GZ8z8aZTngeFa46eMAEvXdg/Yx5NPq/1otFdj02iJm6yXcmiF2FCH9
IlE43UpmACWy5xIU+slWfu5LFtVnxc7p4WyF1ObG+j3lGl0TklY4BrMLkwVBuZXZ
VrAo8TR1RhHU4PXJfdDn1wTDEbR9nifhabCT/a7EFMvJ9IDELvdOxBb+h20tlfwu
Vnj8yOwqGRKkiWH+paicmwUcIQ2BmFvL+Ybhr5zb/fuQi+AQIDAsIZq2xLwhYtcQ
O0MN7jcZdfZOICEIC/bZA/7Rzhq8+4d874Do9umjRRUgE2X4VmWlnCaNQGj8I3Jl
h9TDyqCvo2A0vR89plBS9w+ZSr+9cTrJVUsK+Qyd6IJV4r0SxWsrUtkhP3OfRxt5
dTpTWSj+gHKJMVuf6l9B5N4XXrzW1YJkBA1ZBxjl5OXgUGiKw9jfsJKvFCesEkxl
KpxxewRxomgNvy4n0tCtR3W/e9t0/F2RlBTcW0abZD+a9Y+AZWrP/1/woTPDlo6v
6Aw7KzNCbiO9Dll1cZOZ6DkKrVYiUGR/6i25M7P7AGSs9eAD2caoDdrXuUIrmEoh
pQDQi/ulFFaiKvMLt3cln8KjJwdbWLjXSpHr82NIykAZ8ES3n62Z2OV4JWWvz/zl
S1Eyq2Jp24A3qYgqkCwev1anfPgCcPPv1Z/yA3XnVVUbtrH8l0FkOqc0LoAwlcBE
8sIwNT6F6G5TNjXdUnZRYxCXQUx+/Wwu0y7UgLVTZTlurTDnYN4osypjLRA9xuzz
qdmPoFf9J7K2/aHzxfxghEm7a1nl0dkgunJ0X7PSXd/8GKIc1mVvldkUV9jagqOv
MNe8UXL0Aq+4aHzHW6zOrHM4cm4mTWjGNaFzRjKZeopTV3D+qWVSBLVZ6mG9+i3Z
5wRiKIfU41gd8RSRb8o6g5bnfsE03lkh1C5X18rpP3+02lXdbBn8LAeSXD6439rx
++MVNkw0EkT0yoVsGO4/mFe/eFxJWXaaUB5MYOBeJXh7IWNyJ2+brGE2GgWNDR/1
7SaRc7pQ+x7wlXuLwZBhcfYgUKIb1LbizDvk5mWLn3XRsj6YhRj66yfiCQLrCShh
w22fODDkqA56eymOqG0nxUK3RzcCC7bY2X7Tc5/tb2pk0Ng9PAf7MbH2ZH0nAGWK
b9oKi52hwBw0MvorsM/47rKaO3qweKflq8shil86ixiz9F+okFbJjYlwkWm+jzo3
QOti9xOIHQ0r06WoeR0slaNerpqqKITaan3zmh5ubnsDXdJ2UFlkj+4Jnfuqta8R
zrRgWQB3K/w2DqjyNvdBz1gdczAzWd1j+c8Za0+P3ndhrZT3WsGsV5DpbfO84cCo
/WrAgmSMXsiKM4ERIgpPNPnDR/gHV8xiZs3MX+ftT3+jaBx7E4IuC/xeeQbTgSY2
iRjdH0yzRkukrz1i/xIdUZJsUX8h61qUK4Fg+GS32kPepa6/baXE4bY2Cs9aX8NZ
npqYBMk3nzxoDIqr7LyX7pHkAHgpaMplPQxqlSkXpLusylKXzYv+2GmX4xDSIXQW
pu4n1uq9ivk5xBbQ53EKy/pEH6Nv7TfcxLf3mxMHKx/pZ7y7EWTrJCoxo2HemHhO
T00kS9Ejm9qvlnmfsa5xsubXJZGJKWrwVq1iA8yWQ4vY3kTzbbT7boQDWkYubifN
BFdsGvGjZtfFBa7a8bFSMY14DdNQM8psjM20mHSrcKHVBcC53pvDXY5Vnm4I6rA8
JfqHbVfDy6gaEGK2OQrPMnRnZKB+9eXQb9RMNdjTvJ4fMBWGOegi2BQdAcIhv8dA
Zt++pABjEj/0CP5WqNcQ0erMkjZBi2DCiWFHms6szPYxIgU95TUWnAIGcpfvBtgL
Grh6WO9xWoRjO+5hX1WALXZpl52iH2jQH8dLrDDgvEFQtJnE1K2ECKxfaAubC3Yv
I34ltGlh09m0HuhKijJlsihG+vFeSy7WRtu3ER7F0fdy14cbLJJ+nf4hlPfZqIT6
zUU01SzdFchKrkBu4Z0bJ7T1x+d1/4A+6bGVPNItdy59i+RgGPEMyG/V8mfi9p2x
1mbqUwuB7eo0OfNagkZOsHpvy2U1HEp2ABOeGLYzg9mJMB01CU66UNXQdCDr6L+G
0SwynI+/pOd9eOnD1+OCN1iNFlffFsQ+NHXDe9L/aBstvWF4IPRFsiGEL57Tqt58
6o23od3r89NRWliqVVnR4Gc5W50nssSFr8jDr5C0IpB9pJownUY1oxhZJKJauWSN
ArGSsEbVphNVoY2Z+oRZWhIny1ZZGj9TUrAeC5iugGHrY9jeOR2GDpfTy06UZMab
h08Y/FpUjYjrIW9m3vUk+odI6Aj4bocs/x1omYrtVw3/1Nn2ikkNG2uX4l0G+Yjh
3Slortj8R9sRLfwTPCpu7jEKmcMpRt0FrY2oVQDAEsSRmkFo8xlI30aJQY8YKnDR
uSeCCE/9+OvoFVGFQE58mY1OmRC9oLlO5AgNysuORzlWYCsU1pi0f6I/dehk+my8
YMjgpf0Cbew+aFDdaGpN+i3YQIXCSRcBskLhJryPG3qdi8zXgfNAZRpTP0b6XdSO
KthCFdz45BCKI3xOT9LJHlesHEmVAXTZ7n5W1tFZfZfpj9XbCHm0YyQtD2IUnE+y
AQMkmV9/3HC6JpvG1jEJzhU5n0IdykMRWOKZP/TN7Yy/6GBMQYPJoRIjzreFd3Fb
wEHj6drSFHCVz2UeOYSaDTfY4ih2le1mbqEq3EXW6ibO3EdS4nyGCxjyOec5+No6
AvYtSkz+nGf3GuzrLIGGuwsCuoBG0HO5ySmBUWYNKYWp0nJ90NqMl+XjMKCtDzbS
+GmVNeaXgtFZkZUoVrRhVeQyhmkpGennG9q4GP9btdqUORbwfMRjSGjl+D0Fm5yh
nnxGSc4Ze9mhDkNFIzxpWl/q0gX0M07m3KXh2YvXhht1DWoYpDdFzzrTsBWnb2a2
SIF5cUFndQlJ362nqlQ02j8Ubcm96LsnVGIE/j42/MlJoglPgQ9qcBO/KR9XXK5Y
fLke2GzDzORS6bbzNbdrBBO5GIEwLN3UixZnhbbNGUMJCXWqOu/aSUPtQ1OXdJiF
4Q+2wlZmHjUg0LvJ8bolEIdfDjoH0SH50nt/q463iQ84k461lAk/stX/RQ9AfYaq
M2auVE6SWuG02oOST344uqmJNXOmNo3eVvewRPeoLA9WCGI5qoeSonr9Xu6iidpD
zUmc7SvG44tiJYLSzateJWIN/ly1GF4oU11C9zban1CoFQ3Zl6IFIllw4Lzn3NRp
wMtFG9IChuEaqYvLPSl5VULGoAy2hnuhi99ZeFsi1XfpP7BXRgCQam76Txh1lAMf
TbKW9DNOu0B93rdTwU4UDvUTXo0DoDuhmKcQgo9/AF8qeCrx2PI78qjAfa8lq+tz
dMYRxH76KORjS1PYAXY5sVikSBNijZ9ir6N4VIxQ9MH+oJtbNLfL3kl4vdV87lQH
zWimaH6hktIx9AaZEOglzX7DRH1jcYD/2ynZRo57kTMCEvlDyc1HuKIdmzlvskG/
cQ+sS9JfSx+UN0CB7LBzwdvaOuH20FK2DS2VJRtRcXo3y0HsmtQ9938DJqv1Chx7
0iwbHDsPeAlQxYl0wHOZmm49y37T5Ck7UsYeXRpHJ/L28r/1Y+zp8FxJyt0LzSBK
UsyVvLoIKKThB06Kdto49bSB0TbUC+ViYPUxCEPnPGqV/ooPgg6dAWbbsAuQgXNq
73dINYQE65xpXlkhfWSnYCI4bdlOnUmQMXlRwdBAxarHSxhP+doWOL3RO9e+99nW
FD74gEXUcFDloRpH3oB8dEeN6nVGoVQvEhTzNWNxdVf5Cd1HXXYOOz7165H7+om2
GDnAq+eMIeCGHoTdcpCgTZXzFkJSHkBpwIvehDXi4SEVVOIBJZpmlYEpesuLK/IG
5pQ+3Ly5NJdzmvKHKBDOWvbKf4mjlE5BSimZIDOIQq6wHKAGqbCLetC52I8N3xaG
X2qU3HYUZ2gK3Hs9F8cnkilZWfwhlrvPv+0TaXWa4GUOuhMMT5ei7Xjn1IYkbxhp
eB1h4jJojY1V4lHPheA2u0tj9ZV611/H0jLNX3US5FmRsGbnoSM52ypwepjrP+ZY
FN8Gbfh1qZTxevy508NJsrn7JSzWTMAn0/uDKQ3k/wnA13FouNqypQfAVL+63r41
CoaGJVCspaYXj3aXXSY2o3u5+vQMr52td6Z1INN6U6kHcFrCUV/yEdTeiT4moTYk
7F6LgwFFv/KeX0AKafXzNCO7QBXtIS0Y8Ocg/PPl1jmnjWh58hAmOXfrZzz7UzKH
uX179UuXTG5UN6VWgKwhP4982VVg64CMRRlh4NAFp2lUH4tEzu7pYl650Lkwiey2
vp9eiVtKM2OXWrtEkdGgAHDNX/wvDKOHifU4X1GKiSjyr62jMTjbKw8DYsBZhCPy
oJqC5u4gyCS9Psz7wy2+us17pETiZXO4VkCGgp5vqVj07nSUKjiz3vhFcsoniE36
qLLk434N36a07f+e/mvnKe0btTwXPXkUeb/DqBHpTEqS5y9Crs7tk3Phu8XZiEHC
jhCJriIY+qSIyvQDcX6pHiuC1V4dpNujwcZjsJbDg34hhgwSrVE/JOQBJQ6Bt0wo
7D6Gp/w3V/lqwnYE0FSI+2D2+GUKv+cXIqyFOzoNaymv4oXNp7dfDEcZSnhgeODk
liq/wj1V2F9lRQxzvuRrmPewRMgK2ns66w5NceWTT1iDfY1Kwv+j2PmQQ+bw4dWw
ffqW+MB7bZO4CfRMRY1owMPjtsl3n95Ok3+tVXyo2ANtvUbdwVg+YnzzqBO605kW
u649yQzhnzXzNsjtTCelV1jOivh+/kSsvkTU1NRY7rjh8yH2BpUojuu5/6SNOFgk
hQnKmTWkm4uCPjB+62MhoXKpvFbsIdnl5DV6z4vkLdCdKp7GBWbEYCqZSJYSZiza
gBwwew+iJlLalA2LY5Hnc89HLA6ZBMbPJwjKLB+PQaNqHyd+Q/a/ycVUnN4UXJpR
RUOlft3IXcyuFzbk91O29mPPG551ilmCfIoHk9e4TcVdUVXjcTU2BdQmHpI8gyF4
1KMKSBwTgEOMpeEQWQT+/rj493niiXrFcRblMAG+xPVud2b29Bs2lh2vGy88kvg6
tMdOZviRey+uNePlmf20ozUCCj4QEzgZXmKtYLl/yuVlggghmxpTNWS9GqOYVzuw
xG7KmVsOxRBlf9wHbpOzwbbLtTZXJV0DyOpACUi65woktqx09KQd3ToAqJF9HPjW
EqESZSy+9FdqjZpb1r7ey5WcNNkDcfndcARAXlShG3ahmINRk0I9DMgbs3qMuB8R
o/3s9wa2tPPcKcuslzc2lc2PIn+Ptgg30XAAVd+wA5XsD9Ga2uCYjYv6YUBaW3Km
KbanhCrkOk7K/rCDANZQ1knBarQJNjB2nvWG3CwELbPLdvmzPy7PAIjFtqgx4oqs
BDlW52CDMqG7MCgMrw22hHHcaZOo68FsA0HXQrzaV+z5L35Is7a7T72Cowx6Ycq/
CDeey6aBr/tI2X2ApUCE/mfei4k2oKITke2ZOLL+DRha+BltB/BKdWm4JyMJYTYf
eTgCGIrjtWWHnT792OJyB+4cdth2mtvmKIGq+DCOO0tta9eIKimwksHXLoAhIOVZ
f+bhlTlZd8daQq1vlKx0d1wnsuyNmQWCOWqhlw9wpLvDvSAEZglfdw5raqWmRaoQ
DLDSm2dFp8dMaJhfTeynqx5/59NoYU3P5NjR8ofq+po1c/G8oSLVsUvRd3S1A4wm
T8mpKzYngmN/55lRUDOE/meoomfr/VjNfHN0wcjQ2qwTBVNdUE5aPfY7ovk+539U
RBlvSfdak8r6ZORUfELpMaqeaJQUOoxUP0mLYop8ZSXuLHBWq7FXvwwaaxcGWNcC
w6xXStA8FlhUizEl9CSUI3kpQl/o9b0JlauQofo3Ze5ni+MluANQ5YBBj/k313oi
QtJ5nJkGXOZ0HvhpwjZRBC0HEzA/o2Y9PA3uxBRdwmK3pXAnMdjdG50soURJREDQ
cRMWvRuR3QtGTtbregjyA7YJyKS1KFU7E2xmnITuTp1MmN+fLuTtsD4mPwSRRegn
uD+RWtKS2OwkKSLihVy5rVB4if7NowLob65gMfinAz8wMZ63QqOILxZlMQuNM2kc
VZKid4DzGr6dQK0/h6jMsfzvLUPL9LAtpiwJ9ezOHWtgFl6xPFIlAcpOB0DjYXJa
XiIgUPvRnvTvtr2jxnwAhcHK7vfLdS7EMzlPNxmWTun4T4UrDJqrrFb1PeLpvPW+
m8Xe85uTOju6NJHVtEqkYVvX+EXIbYzY4fYlZ0LfWkp9jE37bVgCk+7SuMluH3y3
94+hY70bLxGiJ2olkMtQxwLBxOYaKGkiVDPK0NjvHU02mc08yyJVW45hguTVTFGP
41biPguYDpgNfgOk0cjz/YSu0Sknm7EyVNez119oZW9Q/qg8oN3RAa+yYQ0hIZzV
qDJqgEpEFeMWCqV/QpyugdovW7v186bsH0hpc8TqSX1rLYNcnVkLr1EfwLIWP71I
fLq3XwoxsV3iZPe/AsmLr2cZtqagsvVV153z6aM8I43NnkeFIKaED1waAKn8Beu4
Na12t/38BpOFn2vzCcBmA8XTgzy0qc/bC7Ih9UU7LdL/5RU6oWlLoqtCQjRonodj
wBjWyrWwUPgQbgg2JUKfSNU6zqKEjbpK4bNlHNIqTmCBLJBNczxaUsuuZ1hUi57W
qfu5QA7AlD5L0SBiymctBOdw7y98CcNgboU5jppP6+MdQ7WxaneLW6aQh0umTZte
hPRITpE05DMeyJXGWai+5nwDJrtcSZ8+yybFsLGxxavpJG2PN/5neYWqeqLuqp05
vagoeDQ2RN+Tdj4leXSFyksgZqi6VjEUhreqERbKRlwlfAEP5OCfyPUCjxFC0+j7
Ig0eVWMtfgcu0mvXoPfb/3zRPQe3GuxH/QvQJGHUT0mXgq4g2gwA2a7a+IWImIyj
QV2aMvswwyLCMfBrCp21rc+5KGRjePMzqjGFyy/kJml+W91mQsLKpCGiFTUv+UI3
R+H+9AoKHENg15jsKYvkwRfwAuMU3TTR2Faz6o5YBmjjUhXj/x6WNKkZDOVTpB8p
chpkeGmHgfbtZQi9d17FxpTXW95SjHUvHm7LI9j08P9c0AlW8Qcv9kp/Dy6wbXMY
oE2jJLB1hVjfwCURfv9Rv2w5LpKPMN65uCzuSMD8HxH9MHJqA24VdNG+YeOKtgwO
B0lbTWT2f/tWC8fVzyhmeF/AWUIHby7vfYko4VwKpAKRBnMmLgw/FEwZaf6HnZRx
6totvME02ovT0E1InekvO0XFiP18bgiXwDo3TJaIeB7hBF3N5u72pU8RqQrL8C8X
izFvPZH75UdXlosKufNcHTZwrRKwR/tlNk70jdvGZM+H8+lFvQAZtak763uVQsvI
7omQybEweX5KQyKkXXpEUrbz5emG1PTP0a/ZmvT4gyAmS4WWCwx5Mh1iqRR2vwqO
jtL4ycB2X1a6Pf49AZA7GPmJ9tN96sms9i6RFtqucZyNblQg/iRH64IW8kNg0b6v
6uJ1m+/9cyxXeC5GarTeW6XQ2tE24q7n7A+ZZl4jceEWKQd8EvO2kicsOkw2Thq5
WO1vF6zqn91qhP5nJNgH+Cc/pwSrDVHzr2XIhFQvo/+3YPggy4/SGyFbf2B9wUVs
tXFgYSFg4yPO0fGQ8AU3/p2ZEMwSmCeAP8TqWbvROzEngJgpEskp7DCVaa4jG9RG
Iiy0nT7iY+m1DEbp/9D4fhv/lamzvKypyBhrMr0NHAmuFOMPPkm4ESlGhVoT2C6h
3KuRzLsKL7fb362ADO6IG+Ba6bFjfcRctkSx4r3K1FrZTwwngJ9CzqvQWI31uHmA
Kz1hk0ODyoUNUHqvft6c6jB9KFR+e0J3OrVsVFF4EZAl+qNYf1T/26ROjaUuhDll
C6m/ZfRUb2Ld3477f8mPvUCi6gpzQq8tYkqum/VdTf5rfoFBu9KPj5XZdXruiOG1
WzOs6rqk9dOYaWX2iClMPu8RbBMx/bMUy0FAPNrNFTH02BOH6I7lmFCL4llbb/9N
LEqA4ukRstW+c27nwDf/kgcVYcmXP7b0aBnt5I67ZlzhwplbuOC0CcexGSan6vBF
w20Oy5dnbH2SHrLIdCLhuTjafbF+49qvsKiXAGhC+OE=
`protect end_protected