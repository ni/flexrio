-- Entity instantiation for None
-- Generated from UserRTL_PXIe7903_Aurora64b66b_Framing_Crcx4_28p0GHz.vhd

None: None
port map (

);
