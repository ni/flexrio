`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 14608 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eislOGByxcl/gRn8UziAa+H
mjgbsd36EQO5Ail/O6Xu+Xx/ROMSlvuBazdeHDaf8f59Nmui9Q5B4mKyD8HkVz3K
Wnv+eGnSPFQTKYMU+RSKVDKr9I1RllMHNWFwa5olf2+Y4kc7mBELTQboyicRQwkQ
RQYNA9aLs4tOwCphd/O25JpnZhOACdugwLrKq1tfezwMB11RYUpjOce0IzaeAcPa
QOmmZpKUaiiiz671so5FueR9jia5txA0ng4mw71vjslIo3vKxG/uGY0nCKT/CBJK
+jebeV33EzpvW2ZIjwUZjW9hLlrtOw93nSQEg84zvQOvfybECfSjEgS6jq5lEoaL
UKhSRAbpKemAOJnEw4Sxl3IJ307rTu6V33KKu+rcnRpm4gSMuWeY1Ot4nEFAA53G
kJvhHgsjJIZM2IPvITkkd4ShhBRy54FpHtM7PZ7LIajjDKShlZqjCJC9gD75HUXG
oYcsHmDT3TXMKVcTsAfIbYZD0Gp5kcNNk3WgYupjVd3yZQZ1M0Vx0MgExDtl0pTw
NXu92FU/7c6oCOa/v/FsxoINgQru/rE10wYJSczvPFm+ML7tlM3NsSxU+7aLAXCX
RNDZ97JU6jihpJcughG84OrhxW9vY4x3GJjxVaKHBcc4OcvHHtPfS3WJbj9cMgAy
wKCHeLuNWIGaKg6QJJITIZj9BKydJPBSZQZyyS1QoE+Nung2DVNY4yyjIPFYUW54
3K40JdB49xn+B6+aU8k/7hxMpPZOmn0PRMfO/HJUSmibHtKRyRSX1rsBw65eDl6V
r1gH8326CndGykjfglDOHj4f6AbvOAkY/94fPqXM/yVtbnl7gh5oqNG4jvAvtjnl
3x/mrn3Chk/VzKFhRBPReGnASFPixQqpZKdwmluI8DrXby0N0UjicIqX1L9zO9BV
QqgjyVoCyPqJkCz+2jiIHuJyIk2+1cyW8AOUeGjGxHibREbGFsURRHz/1AAfS1oW
57wPLjgs+CaM9LkQV2RnySsb6VKJXegleuSIV+dnTBWJpDR8EWC8uOM9o9mCRKca
6KvWtCCffhdaogOl+bskaWSKh+tptMVSNeobO2tp7W9157xhYJdf1xs9N2BT1jfe
OZ1iWKCGCAX/quOiwU9W89sFcsuqm2xQeW9FaR6+b38Id3uLiSfvQ/zzlB8r94wW
DAwmlDJOCMi4KWlwntAHRRE2ad5J/5aetcaRZ4dj1k94pG76i+f8TjRIJ3I9gkXg
C1bqG7WFIH8a6mhOlKTVELEEkc/6uJPVjoEjEcUgVa5wRKTAMDoCeb78CIjdxFZA
UEeWPYkMcHyda6Oe6oAL54dLcoV4b+OcUy67L0f9UPLKnyggJEn+8RiIPW5zEjhU
dJcQo1JbKnSBtmyL/ncbsegb0kNwlYxWNUOlwyVMeP9gclfUyKd0Q4NhsfjVcG3R
IjEBnMb4wv1REvQqY7Q/eZpyr2blVtpfcHzBSBEN4JYHD1RhqbuQuXu3S+rm4Eg0
9pg4lVSJWtxeA05Y9RYzAp2GmD3L9ZJ9KWkd7ycjaGumjNBSjLEwNcMOqLfZnEi/
ounu8GaYyWiwgCQzFl1/KUNrpUuTgLherOdjOuGd8fVemG2D2nEks4yjLA/Q9npS
XYflsUg9DjcH81R/orp9gsRVaAh0ZYZW7QQQuh3jrbzLIBp6n6R8S2NRpJXU+Ox2
/gTbLsTkbSqakSr2icUTv/+rnW1UBG9o2HbmOuPav5nbqc7rgQEJ6AcHXHQK1aBJ
sKT2Q9Ct/TPjlgEeMvGlUQNCQibvOixVV4M/sN/TXWkJV0/rC8ef3N52IpYVKFsH
DUaHumhLtsN4X+MAwFiSVS0hbSc7hZoTPiML2LHLM8FWwM5bE/JIbcfU9UGRP01e
UtNTv+V/5TxVsBbVZuLyuURjekVxSVWC95AupPLHXKC+6c9V3g5smY2XlqsErEbp
ZK3yhB9jcVhhRzXR99xp3ZfLu5f5HGvZcprIsvYZbXTzDfa/QmMscUqHrX3k/VWi
v+UDf5+qv99Iv0YV0W93LUSp2bXHNXRokhfaBTjFoRtEMtbJdx3VZb/THgQw5KEc
0veJDJGz8/sSCZS5/P4hwdmAesJD9dmKZz9mQLgKL0JMy6iMIXhGcf0By7G5c7Ir
pT6KSVCiQ2Dd5qwn74jKe6HIqLkSlGg9ZmIowPDzsYx37ZIP5HKE8MmAeGvNtptr
eYcnx3Az6ovAAgNtJlJx3KXSWiTztrxi9jbRP0LPHyHbzeyCE9B5h9eX+jeYgyGB
cA1aNZ51s6hqrUhH6tFimQUYQNpeeD2ugZK3Pcv/jnqQ9EdjH3Qk0mPLm/vxy4AK
bdG+qVUbUOuf69GyXiXGSHd0MTHXPOJy6jTPQi8msSlU18bDwrSohjFQGz7UfIej
sp1PybmnBcTC8e9MONmL5otkId2pol/kMY/VyUif5O5D+gBMQxlwvYkFjiZcxoVu
x+9xudAxZlLZVISDFp172+X8egaGY4+6n/zwBZNgTcIzIA38uyWARbKX8CRZBSlK
YmWvqOAYieGO+syqY8yctS/dxic+F11Dge2Ym1A6aIZySx/z4z4odKlgDEJ9DNZd
7Mh8J7vIt+CDTcxgtL4WvvdGgFVoRF9El3pKWNB7zWFx7jcUKquFzgrai8C18CiI
BkiSMPFEpivtWjFEylkgeam019O3vT6dqtg1i99p4yfu3ks2aa/CvQ6Q3lrjoMv0
Su1niDkFVQIgkzdRzLolCsQgAhABliXtK8MaCweXF4R/xiC083kZFTc9v2SN5JLE
aLqslvoVPG8JNoC7T5Cv3LaujDOj7tG5BDDRgzFLFPF9BqidCCncIsM499Vnr8NL
3QfjxhMC0gs/hVJ5gFB4dJkFnr5fEL2lSsFYDR+H0JdF+62KTID/9aaLAeHYiPKf
NlV5iTG4QF0Dt3J6eHV1voWKS5HQQ6AAGctGDHYCCxTjEUxduPeGTEbLtjzU9VC9
OWTrlBMP1XUWG665s7A+hDfff5reZ9v2Yi59qqbf0kzT8hHAqj64Q477v3+ga6Ym
4jW1oOjWkX5FBTPazQXnXAwmFUSvDbU+hl8GRAXiqXPI0g+TIKoHhjLHJWwMNbq5
K8uhiF7KHmCakh6+LNXAagnqNdNGN2d8wHMczPGiGficADEWNFMVCrWjoXj1X1jG
PowpYkFpugt72tKKKqbs9FwTuOuaBaeuyNa/gnfgQ79cM2twKHWtyqxtOqTY4OyD
k2w4ZSm1ti2AkR10TqKq9DjS0Nb4lzjOMnNLAeiCeXJy5eoLhoP13xyWiwpWzQuM
gtN+C6CWKG6jACPJMHcJOTGX29q8f7nMhm2GiJzOOQRJHA4zQ8nQMYAmjBTsyCzG
0C12wwXeyDZUJJ9E7UeG9ozC+PtPGmNB05OXt4fza5h4yU1qrByfGU+h2jsE8iz4
HGcmiM+S1jELYOqD8k707lwoj2QQa5QZgooBduGaVIbJOIPVeS4rPS75huTOOGtt
LXPu28wEi0focSUGwFchl3bvj2KedUh1238sHnrujbhLWj99ken2wzoc+XJlGWbz
guCIOGTU2ORJYSM77hcEjgF7HJ3vBaVReXQXS2QWFz9Z0/0uFEejpy3RpKE1Zh0o
cn9i+21op0wor/Aa3r7pxWBn+yuoqiBy5+GQv5IGq1a6gGz+tGradh7Fvzz0gqgW
Z3+Bo4z+wNmOc5p6xANX8Cmpo+zf//v+szsx3Cx8HZ/hHNK81EUpveue4xPvWuEW
oGZZ+kL3U3TWqtxFPlcSFL2Un7kxdycybF7IkrWQnmzLVjD82yZEBn4ahanPMgTY
nn2eZjPOBtwo/m6GCb5qeniNb+y/CXu/ZSp4/MZ2FEAQFwLB//Y0oXnWL3ouUo+D
Aa62ZP0qal0yIRWevXkD2pFMPnZj5yIi8w468exd5RQpVMSQsRhwP7SOM4VarXUy
IrzZdFkczIIPZXkVmxv7EdHEkSnNjuAOiDL4p7v7NzYGHN1SFHwFJWmF/mlXtg/f
rZQkS8hodRutv66Gbn1uRux4IBDvpgZafjWdTxcozSCEgDQCCtaxWiHM6broamQ9
MetgQIYyqlPp97YcA66PyB9DJFvlFDtf2ygW4PJFlrSrmn1BRZtQ97gZY2wkat2F
PEV5ymvBjK3cgs4ZODL2H4x7jnnLJWGGoj9HUa7qVcoVv0BhaHG3FrSFILA9kro3
MUeeoJbYLMefFb5N56elgESndo4i/g4r8sWe2qp4RJrJBC7ouNllBic4zIz+CM2S
d7lb8chC30jgL/psKczFIdMI9z0ni7iKmFEpUIOOWgtKVAGQj1OnOvFXyfjqzPPb
Y5JDe+RBznWKTehs6hun8aXjAAdD0bwH41BrR7zZyk1n8DwP1DUaaxftfc5oZ/4o
NkC4tLG0M2gZe+s6o9FxCB59m4V5nMUFTFJ5C6wD5rPXrpZNDOq3xX6t//u/aYaK
UtN5sYFAXzWfw4IVifG4kjK/8W2CRaeB/BSYTXlX96cAzDuNj/S8t59NBU843nhU
KTyx7SzyTM1szFjIniHutlsEivuRqLgsd1leIm4UBeAw/EU47jQBCmFq1s/hVxoE
11SJmRSyg+BzTjTtcIKzjg9S11kk7fg/zLkzb7libkfJbMEeIrTa/Scwke30ZgLw
txZeS/p1Q9Sy3M9l9ALGeBUgTqDuYYOZcI+eKG7zfVhRyGLmE3vnCNzWfgz5OUKr
Qp0Sp85T/a63+g6pksv+OLzYIN1hgKPcLLFbcDxl9BY/DQbs/P7lOFj9v6DzwSCN
cb8o6PedotZen2xd6EnMIpCji7VuoCuFaeH8GA9E4QmItWjzpvcpROPuTaR4tl6a
dhnI03BG4g8v/UnhK5mWgSez2Yq6Ku6As+V/90eA8ceI3aiEZkcT/Tclu7WdwJP0
Q35YgDHkmXF8yudGeTeYDlrnqkBqDr6zVEbHuqX3kbOIUCKcVs9hbOIoVf5JtDpt
trsAOUoZOCk6My+fzwlawZSGI1Rd4cCrWOPPM/8op0qOPmRaBhzczEmp52x8gHvF
IYLbhWdOF+1dcSluRzEzTKHm6FyEIjWug7s4HQgkQOgyYEm000UpMn5lK1sw/GRm
2Gv9P7VrZNdpWUBC2AUtConspVDOW2nqwjUEBAPCZ2UETjY+YRjSivFYETjlKz3u
NOg8+MyUsffm2CALXT8nLFp2aY+sX8W6S47Ao/rdWwBUZXIWtL28oktfqLDu0EdW
y33lsn/6dJ3rrM3hm3SCAkYX13Ns2BDTH/Tth3rNmGAoGXZueockKMKKGvvjexf2
e2fbdQkeHgEuSpGVfoF/IdPjGKaKfx0ruse7HZTS+AOhkDZnOBQcYqQSZtSJwnUO
8iVtFCTPZNpkPnne45KVGqboIr1FL2Q2iI1hvSLSjItdLvrvyGEc6zAmWfmutIX1
IB7CNm2erTMOAoLp8pW3EdIqDP9JnOWry5+VI6UfZtI2H9slFaCWKhoSlqbdmqho
yGQk/lvLY/4MDPML78BoT42xdf5xmUT0/woOGalV9PaCSweOCmk26RmMaAYztlHo
Is/QL+6VTJ/rAf5IApMwCPifEeU6EsTfeIWE5vhL3yLt/X8uMwzKe0MqBWQNkGPn
7G2ltlF4waFYt97lX3NaH7nJvLa/D1B+6moZOFFmeReS1LeH46dIUg7XbusmeV9m
vf+hxkn+zBHf217uoKclkt+kaWPxHyIkroWHUZ7px0ZDt89u96jBGBpE8x5KHCNa
DrPEiuBAVLdquLv1OYxLVCtL7pNiPFXwICinYrNXn3Yn6FGl9FWwxzW7IeiCrv6m
wi33ibmKEUWmEoSWPK/wOD0GNyFAcIyreNxLmShfcYLN6eFO63QMeYRKXJ08CePz
lM8dD/XQM2ZEkJsbyfx9jRpV9Syt3hLCILPy46lGq284yuZrMoSSAuDim2Fm4f3W
ZqINSWdzf01eNOHgGDqH81Lo4k8Lem7kyJTusosGl9a1CZIBhc9vqoP+7P5sf9tI
IXVHXybmdGok1NJmqqDxQf80RHnBo9VaFRS0LysWr3Zt4m2QLtAPGdjCHpM+5Gyh
kftNSjNzBmesEg1JrIRS+xTPKD+l8T9y6AeGnvbYaXom+8yUG4OHJGsWSIUvUblV
k+opLejzvN9bmadBMl/vmByYSVDCJD1/OCx6MzThAmOZe97udTqpmaxmdvRg1Xds
xWALSgg+g3EXAPhissnFJpXL69nVHAHfgO5x5h/F6ruDt/uT3ZgAABi24EhXtrhY
nZtxgAWZWUFlhqXxAf3IGwqUZIFAyxQ3vs2Z41gWYLeCcnsIRbrQgVHPp5z+RK7O
pa56RYhwFkfwmf+rYQvThqCUxP1MiU7GGz5wrmAaEfDUnUYXRal0jB6U5jBCuNOy
UcItwKa4u5MjlUTptgOshUAHXy2IRLuej4jUfX9F6vRSLVRAF9o7lcfP2JFirswk
F+gsDrNC61AdSkFq34xzyG4HKgjn7vafevfAzmySgGTk29G1aAMZ3kHA8P5oTXg6
ndtbpicYYWecsiwUTyKZnrME7r9AeiggzfI3WWjw0SA1O6wt95u6WZBdED4LisoI
b4EBfnUgJbNbzqMe9v6PgmQIOdTFsD/zF7NUvlOMfLA9Uu2DzwdmGTeBSwITpzHl
0bFERw/m/QclgQgPhICxPoJf1R9cXoqJ9XTbwR6vYXRSYUuBlJ0T82Ct6Kp7wnu0
vliifm7mLp3wwncvfoO9SoDX8bhUrj75z4en5ik5V6+Vz6VlvIUxRG8qniUeTnKK
k2y5CvjHwr4nRIyX8zpJZpSJLezN3e2JDBPU2aKubhH0YTQHvPkb19Z+jMQcbhga
v4yttz+4l0qseZUNOyBsYM9iPetDakHza5rZLN4pbeJOy+0AK09ElUdTFAuiGY6h
1URUIeV26QHnK0BUe6LJj+2PHkKFjbRlAQJlR98ULBy7u1rE1GB+m3UNMscGkHJv
BReyVWesa7WotaN3X3AKEA+SqIzKzGVNwg8rwKfCxmc4W/GBy1lEvpXYQNltS/1a
cY4CT+DDA8c0B7XMVWUShTkGGebLyLA12AdlXWS9ktSBlQxWWxQ2pJISTd5jntpg
towGG9lYD7nU6ExISO5pbOCN8YA5vJpY6TYB6n1QQ/zMlpKEBG6S7VwELx11rXHX
b+Gnfwlp854S7ynBV7OBhloaeBcwgF8ENzvZYo+Hrppb/izaEbriRNzp8zVIvn1u
jQFlyuOCjPrhH8mj97M4YF9JRd+IO3TfL30IhEXT/mFCIdbhm9urelvFjF85Zf8o
JnaOE1Wt37+dOTc5dx8+k+bvxqK8KOb8wKiyCYs28cDajXrqv0EZOlVYuJn8jxjW
/L7ivpgQ7VW01x/cnAyeuFEUSxqCcO+f4oCbeUVo9EnsFoxA8fHqNHAao4i6HowG
j8KiEoFAw7riBNhmyzFH2Y4mRPhCTLrG9Du3tK+4zySVe5fkZdLEf6DHEX3PaBID
U+fJYH76b6P7CsoJa9pmMfFn09sBEK/w+JhlPzEoaxgzwWik2d1QpaE0uRVAZ1y7
uuT/hpUM0mUKsXZJD4qXBaf59WnhUlB0SWCX0l7caShokE0cKgcNlDyUujfqBFBl
WBpPT9wEJmrEdbjvJ0kPOsLDsSM6LSq7yXGRHvplRksOLW1cqSzWOCLyOzg9xdCr
phiqKIeHm9LyegTMloJ3STsEkiUz7qAsJajSaR961LDZikZLqnpPD1i8thprVMk4
op3Cj4rli9Sg6zLp6SHL6IKzzNe6uDAIzVnaZgo7G0cyKNaClEkQp5JtTMsptj7B
skP409ASGfbs3rxziZZIijpt/OOt60EP0U82C4bXQlZzQhgQLEfZ53JnhjMz5dr5
Kn146s2qt3ZCTXj3wfziIjrpxli4pghiP7wyNNZzymPaZE1iFc3/ErO45Jls/OxP
BcKOw2+gHW9FP5/Dp1RCuizWg+nMFh3eaYQKbJ1dy3mHGxlcCLdC0rM6V/XkGw3o
ZinLFyY+BGnH8QdPVpU+Y2tu6LAEkDwY+z/aeC3bzW7A3FE0VQU/zQgI5fW/y4AC
V4oz/dQtvHvcvQqMDry0OzJkfjcG6ZZVYsI7c4Xc/YEZxYlyBlmlLmLeIj8kRTUM
QB5tdVik2QDzT+bfdIig/2HFYbROmXi0t+AFEJr/E8gN3fKsHxUfByHbkTpBrY9P
XrbhTeFIi2KfaqO1brxfPr6MKfR1MuEKAyZJROrZMQHwktHN9WC6TnZnFqkXDbDW
g4zbTP3KeWTIxa6VT/cbZ2o1/7roa2XeVYytOBQd/ILkcipDltUGTLqbwsVRpaK+
YP8ar8yreeNyljZ0MfSjWs7BGLQdky0EGvDSIMVdjYEYe3KLyaNbsCiuakMgel0j
fbINsKDHR90k4vi4mlRTmR8xH3WcZ9IaBHaBKSdqiAcrHnSqXcYS4KptW+OPmoKn
8sXtrR4mRyrfTGXoZ2K+SNccf0ylOq0hhlxXYOPiU3qLx69OsXfEVL6svFRQZObT
oXXsatbD7Yy1zcubVsCHaNAzkXNeJLQBlli7PrqB+9wvhdMQDTUKdsm6PM6NuZ4e
U4HAb0IY6WGc3FfpJnzYKVBtST3CJeT/9M+miMzXTQa24XDhLepq7TShPscPgYVB
n3CJnEFEkKqo8buL+COE2KOsUV7ipC45U0OricGh/7p3UUN/syArj0hGrV9Je8gP
H0MYhWqMq+Z6Woo1W4gHyFPrFzUqS+JS0cRq3+/qEmki/zgYrQMWDQ7aLj1fN3Ng
fNrfHrJF/9ysgm5qoFKuYAG/Y/M7/AX+k2EmuoKAW2doi126kKXlmZf3jSgEbtSG
iFMguF/w5w5IJq20/sfNSpwOfkGnyulNUUVRCG3FSTGzbm6IzoFS2vmVGoc3Eh2C
Ac/pQ5f/7c8UHXdngvO0HjH9+iLTIn4+8/wGTTU3b5epbw3SK4wd+ixB0l0xR5bW
EJqqSEvDRNeKx+klHAcFJbZTF33j6JPZJ75Of/YMz79XqqZwyRaRzNHpW+3UxH96
TMGglQJvg+FU28Xjgzm2jAiO6lJS/o/fv8LM1tQ4gavMm6OmjbRejkETfwlwlwIq
mL310LUgYBqhoUeO9HTT4iv3p0Vtq42/xojGq4ZniSo4uxDjdIYsHgl8BXuPCBpI
PtXNw5n6BUEOjUlMRqGVkmq58YCcsnan8iRszVSnSrBbh5rdeptrqQp1xkrANx10
gcc5XJjUvlOCnvu+z+wzc5BXqyayYfFtXU90F8EHJCA4AXct6KjVDEHuY0fKjiFM
yq39BRM7VSUlW/AUUPM2DkOnln0T5bo/TXs8sVJa4/KD1BdJ6WnY7wFOzghydlyM
wjZvvTA97WGQ8YEv+YG7mGXRltqSKT24YLD0NHojqCd8UlvwTPfT1cWLSgsgSfy2
Bzr5VjQ1P+oRlr3GnzkC/JES+mKtnmWvLE3E2xfJbOUGJqc/H0EjWu+OMrBqbUDm
+dh2m/SzORE+swDXt9gpyQkNWomcQlcWCCxeaaGkiHwSBdnREnf/NnCxOLl5URhV
Ik64wbx2YYEgEyrNk0PGE6dXeEC70OvO4lcG2Xq6lqoYASIxHbVOiGoq8dCrrFnp
c7J1YX56YQmi8lpbFwJr+FfmBCzDSP9EmsEw0mETyx5/XVgfZjx4OyB/1Rx7jGrV
HUphaKmXPJvCHu0iRqbpA/YMYhNZDHxzelHrd7d/0KT6L2u37bzZPqONZWiDkEwb
QjIAWivqkyvDzPMycNE7TZa8wMs1ZBmaXRox/cFjbsRksdUEs5vOQ429BHlgShH8
KN/+B4dVB1hX5GyGL7zFV3e/sQBigVU9+lJCnwyed7WNYgmEkxEUkuImIZK8fCC7
rtyZpj1sxw74fAF77ROrY0UJey+wvmac7NfngvPl4QdaCfqfjPx4HRjb/WiiMlNQ
cjPK5g3VXRk8l/ohoBO+npRUzoWWWGBzCUy/yD2kpK+g1/JqnQvBvhO8gcFqLN2f
05Xjc3lYQyf9wsqksfTG0Wry8ancUkNj/1fZsRYcyacf4+0OCBQsOxBq7jv52rX2
G5gl8wPAd1tfWLpSJwv0Ttw614Ri6SAGkF7sLlS6mJY31l6kB6BWfrxVU0x7kOut
bQ4YfNJXQTYeuQ3MyZ2YAznhOvEukuNbslZiv65W5pcflKS19prsHog9dqbRjsyA
IaTeYe/LHHMPbC1AJ3MFCnAWqNqCnQQtl8VUtklwqNMDzET98XbcYmgomF2F3zX2
LBORxt0UC4IkJzvQX0mHCLtnfv7rpFAifJjnOaIMBqqNmSLey5IpQ+T3cJkyyr3z
eCn8kO/vCr9p01aMlQk9acJ+c8XbIRx9abW7QIEm/eG1ObWEgU88Iafegi8kCVHG
4SY8aXaYF2yr3NCOxlZLcsPF2tDuIjOfkalFi0ls/jsapoJp0QNr20kaCeApbVZg
NFhkxHnVbm2xYTkCBGq+rxvSAScTPITroU+CbSS30JDjV/wOFXXM+U323JMMhoD0
uCwc1BDZj3FUFQ5Yrkq69OtdmJZQmSMoP3mnGudrtImqvAWhHfYT2psMqNte94HB
IvZuSXfMk3y7/vfQtlawWJS7wFRkzH1vZp6xyQ2Xm8QLmw5XJI73KkTMe2SUL0h1
wV2TrjUjkYQRMnEoB2H1cF3RZylxRHI0EDqIAIvpeF/K3EpFgPjbl+jq+FPYB/wD
7T/08Yzb0t1Vz31g3Yd29EGyF06wXdXZKidm9N2n8h3Oh7eoYJe3kF23BFyvGcMd
c9b7tbD9WrTAHxOwZkXQVVSHECwSWGkVE+RoLp64PpCsuQpPQvpDfC1X+pr/2hIq
6ghM+Ibv9kSVquqLapPpvbN2Q2TKOtXohwSFttjHfUGsbo+VM88WSnu5Dpt2qMVd
f8y+bF/UG4CVDPIUDTMgfG9nQrHgyhM/pfY4ck6f9FbPleLDY11TYSANUUNG1e94
PYjuOGLv65CRuoirBtxIKZm9dxWIYlxQADieBoUMxBkYAnz2KtPbQjteK1EcjiZl
8MAvIPE776PsKgwHR9+eC9eS7ovQ9JAOwB0AEayqb5o6khPvWWTMYf/SBt2mymNj
Hmbmhfq0LYWGmxTb7hQfv/1Cz4aZ+7KpHUbgrrxEHXV8fUksN9TFDqhG8tO3UsGx
KEgcBhHeaAZglAOyvnM3L99/0E/+hR3cC7+oCrIAu6udps6XWkYk3HusbOJ/FoHH
lPdhPNv1qH7QeMKnQcNyESkbsgEk2zO6cM1zaAz2Xsp84c/CB5KHG3Zb7lobOa0T
Znh9mqo6fq43Lk5M9In8TadUgZ/LyMrAh2jYl1goMF59lDn1F/7rOIONcO747GBn
9gozGwFO3sljK9BhC5jDKTcWZ4OoRI7Bk5TkPjiG7wvLDlxI4qGVl+J3bhPr0j4C
vBaKxAXdsjw5QUiFHuB2FCnRlsu7JmNkrh/kYFfXJEottpoopl618lfkGTHaZnaX
7wuxo727YQ/CHRUaVMgadH19KqohzECTyLyqPtxrnkYnAh7P7qwz5PR8Gtk79qCc
YTwV7Rlr+a6DBxKHvAc5pMVWJ4WSNHqOFqn8AlX4eRZLlcbfWXssegJoh3fnmoLh
DmKr2sOsgZrkN6UW1RhrpLuenqLkBM/1BvuoAh37nw9MuLiCMpvtYroCkjahnamT
MMOOfG944bCejG6hjYCF21OU026TmQ7qTMy0Ilqf5fKne7xvCPQ5NiuBJWjRAFSd
xhtKaayLl4rAJVdbdGKOXUOeD8Mn99K9VYaLk9rhX1KE9v3Bp/ALfff0xwPbBIBB
vI0kd4noM3auea7k1b39xNAe4H/XNKseJXsE5fmYQ2fvaLI+1IjNVzLKamQZH8VH
J5BH7wB4eHVFgM4uEHlv30zFLvF61SrrRuJBu6/K/dXl5LXHqM3432pI93OGCQog
8YQwOYptXYRc4jdZmL7/oBNEDv3H4YDKJWSnT4C0pL42F8UyL2HENDAjZfaNONV9
zSPdTWkOY4716XiWSfazxVUyerjeqDXxlc7YS4Q8oyIH7LtzV9eMkWN/MW7AUfin
6/bKIz0VURxV6QdyafUdom1twI+bN1Fcq0LC7Wqb28xN5g2aMRU751EnzErX5Bed
qIBnWkQVIdgyLKOY/+51VSWkJOiia/+KYWGp2Paq+bdxJDsw5U0ZDsMfmzCveXAk
953htO8GOiHchUKfsNwsxwcrYhmGzJEF/RjmvkEf7Uz/bDbMsKcI8gv7C1hp0NF1
8SyKTcZWqz8PeHhRzkMAVW4knqXksH+zqqacK24AG67t/+mu0yUUP+5mT+fdY9Y/
c99MuZO9dww0OgMowt8hfSmt4/p+lzTu6z7nC5O4TcLgqIhUaM2p1hsw5Tv/Ckpq
AoJkFtqjIHtmTd1jFL4ARRDO7BWROn8tZ7LnCVHsLoQ8HFQjWLVhBbVIKrmFz3p3
kyJHNKPYR2+VgeLbAe8C0aJw72nMunIDSHQ/BhCRhsPuh4ygbqBg2aJ8iKBMmgwd
Vdf9/bJ2EEoImIkLMB3cFkQKeaJGJUXISBjKj32yEcPLIEz+VoGDwUD4SFK+zQbP
EmazOxB7WkTU/yUriZHOUhxIdh0mx9bZSSFFoP5iMTflj10+u1WMxXSpoAYMSVTF
04srNIHKzlHhHOTLS5Gwtq6IAzrBMIA01EC0UsNqY/ZoZog+fW4mBTm///35Eu3I
B4s3K22fRTDGop7//YjjL03thpixX/dc8Lp8MHOCHJVg7ZErVjc+N01P3acgsLIG
a0AezmyT+lwjPWKR/pwOvrkdtg47QjHHUCr0nyTCumBGUfbPINJw08qx9uP4K/ry
RqQKQUOc8Ym8qeE2na3UsnGYY/v0KyEEdPpW+FxZFX3HVPO8qR1CtviV78FYNB9j
rhaQA6b3iJwz9Al9GoFIgTzEEDuXyp5WSomipWPLN9ygjefca2VMWIDhuq/1HYWE
ulVmLkjeud9rf8bnC2N8llFBalX3hPpWdOsWPMoVSf+dTa8P/q+ECnzsTQ1S3UTL
UXk8+uv5T2GOO8NQ9i7QndDB7lgTgLjHFSKWz/TONEHLOqku4dxXU/JTXpYgKzPw
sluE2dHvQ+62SdlyDj0EDkKVwOKRMVfSiav1p1GTnLJiXcv05Oq8vyhZ8dPT6rj0
CRaEyJU2elO6jLGtzg/LcqD6/grc97N/dmDBwVlc2IuCivEwtaq0VbIRQQS7gVu2
lvTom47FKYwrVkL810/F/k/SeFrZc2HVSsU3p7Cbg76qe+gRTaQbU1S/Fiiz1X7b
NtKevVk+aWaDLYVgVbngwwdcZ6VS22+TlOAg05st1jrk2DZYOnMc8SaEVNc7ml7C
Ji5Mx2Gnx10R2x7vvxRehh8zUN0sZBE40lgtzFpxk0s8qW4FfWcMssMOhGRclTKx
/t8oCm6p2TuH0syafcmkdgSsYeOtRe5bc0bj7LhglPB/7dAeDykLfDQ0NRjfjfXo
Jbr4v8eqdsDyfSeMNFJ54MPTaahfVS7NcAKULWSdAjgg3RVl7tt3EDoH08y9BKK3
C8YRBcQ4K7enEzzn+dxCc9FXnVy063AAS7DGKrookM4BQc0JCWekD/0eleTb/LeT
VALtAOhQGKkCZG8vOQt27o9G6I9QUkL4CDodCoMOsFaVkgac935l03mp+a7h+QKO
Js5loeAVlMsLcwjNJ7+V5s4wg0ZKTQHJCi7Klk1pkl3c3EBrHr07uWwxsoOMkr2d
hypnZulGjl/2kybZdmg05NtVMZgF2DhhkEPHsNKinMfmwokm9NHyhTJFYSSdEUMZ
DU/hGf/a4QwfzdMt5KKy4jnQg8f0bbdj3yWPpaiWHR31PPNWZ0V6f02eK/hvzQyr
N1t8xn+VNzlVpWqQXMHK5HzB5AEGGDjZ6lky8ipZNUh5XDfQkRoAv9h3yBzU7Bgv
bWmsUelTjGJbZhzj6S28ODM7spU1jdZyi16N9kn9rZ8xXxZfZ7o95i26WXkP8tlq
09EdZVUWjA6g1D0xFvMOFONtMtlODxQt6Bg8AyUXWXxqnvOJD3VBMZMDm8WWcOLf
/gZepwunwGknID4kNg+qMKc+MEzNf+psbV+XWdVhePOGyEKLNJJjO3OBHk3lnXX0
BSWxdio9qvmYFpcsYUrLJD5Rk6t5ji24yzDFQFBBqFCD3hrKRz6iCHaSC8mdsS4I
HbvtRhD8yC+D8NXwmWa1BcjuUCRzAwxPP7YgFlWzrsVp+s3XPlAOExcKgSuHqdaO
5p+DFAxTgznWbHK1tDnFZf/He7NdAQolpOwNKI+UtFY62aD6+DOzlIwWuRcG9ewI
mUptZFBqpvx5ZEqFHW2qRvSv3bUa3+Y48XtBBj/SYShri2EpbRvvYji4pNvE0no/
465y22Q4ACQ3E5PTxNigQvFlqB9aWsZIHlTdnKPATHQSaA21/WrxMSPKIL2CwDRf
UVNWMBO8QTjGNWi3djKKGZWzjEXJ/GRQLVrDsPRW0Cu2Wzuz3hGPdYLmrjkn7KvI
fCTltVxjsMs85rLEX5Dpt3vrvdZyKaBFinjCQvdqIEPra4jWxo55WGpWG2RAO88w
ToCi6/LuH4MF5ror9q4vt+OjJ6k4DPE1mKhtZsI2YOupQUUwhHD56/lOTaM3IoLd
cfXSf4EQi4xsofXYCfh06OrU+jWPmNGudn4Zy6AwXtz9qnD4MG+d6VU/3vDnqgiT
ZJEk+Q/P14vGTvTwFTrOmHqtrvFa3RtimUP+oZXjjld5YKlE737ydVMhUCOnCkAd
o3/C5QKzq3e4+u22NymQ2BHnD1y+McL9vNDb84eMbbF9D/mOvFCs791OmbhnTLYz
WW0Jh24Zdcvx4eJQyAoZ7To8UaOpyjBxq5EJqxPksL0NZNrBPtrUqN9I4DdgGHjo
dd+ZrD2LED/qCSydZDi56/Crgv7xt/WEKM48I4XggYfxpkoHYIiDHzq75Nz5V1cp
61miY0YJpSsslnqML0uoVWy4rUksIjqbYD2V6kx6dTECqAS+cvWQlnVG0BkxPGJy
grqZtu7VTdj+7ZsGvFlOkliUpLG+IxiknyvM1qG42YpDZJfTsm982Q8GsacvS8SC
6+TUs0+IThfNjs0UgxRpuTIsIi0IRkcL8WnOo6M7aFYvROgqJtpZCMBe5MTwWqSU
C/ILpQaRsGAV6wil3NpYgUiFxeeg0/O7VUML7/V+dfXvGkoCPgFatIEkWWPfblrD
krxcVTM2ubu3gFi+J+nYj+O4sR0SLiCLmB+ZqfR+gXTHMDwkYdHJ+bQWihGlTpde
DyZIzWurbn8l73a4URhu3R7aguLbJukIxaScwejl0mVnoEpO5YvYhAJSjU2TmYIf
7VvliLn6ac6hsxycNMYThdC6rJoZM2vsVvoYNH4Fu7sAwK4JdA2dJBqIIVo7NqE2
rIVJmDCAmTfgJvIq69PtqODbD0jbqQycXGL+4UJJbJwyIWvKgS/KFv64d6+Elkom
IAGbIIvGwAZ5VOsLn+EM/Ikqd4YFLOBJmIxLJFCDerkJH2rftcajxFOoN9vuV1C7
wMmpcdxdquWBvIdRncswz2YSI998FGMp//JU48QFEtyTuuLCpDVFEUK9Vbt0Vfrz
ytI12c8sSTTmrMvNJAEH1RJa/cXaSsOTtPlIjHdJGpfjkrT8PIjfMdOjt3/I0+Jk
7O0OQb7JlblPRy9fRScfl6vQQKEyFznCuznDDwkRXuASG0M3F+aBcIV6z+ENraYK
kcNqqbzKpKvcUMiB0Su0euR82WszsRBCFg36Qdo0C8gdkIWnL+6Moo1aG06wkJwY
XZd89ry91qgSAnukoWIWw6iWhSsAKmIYden00qtKwJaxPXytUv4VmJ6nUVRk/agp
9mmeXuR83eaCMfY9Aw7lBe13ulYFxLD+8woz94M/g1wZeHKXjo241F3Ct/E4+DJK
8T4Hcd0eqDJIrT8EXIIVO59BdtFRtjazv8YE8QWOpnM2RCdWg7vmMEW5b8WIAWjs
qRdD7YNRf0yA+K+Vya+6iMtGDRs8avCtboqAQyoJu85zcmKSXIMCdjaFwV8pxYJB
of2Xn/fPa/ARZJtHME/phvQ7TR0iDKtU7mWbYaFVTIDUun/yeTb/pZoSd4CCt2wT
HdVpi2xkPfW99AJn4jqlOERGBlkGkEMH5EN7qckeL+5iHPHcRy9VXg5VsBGWwIa2
dKzMdGM94cWsPtp47CyubkTkPy1Ptwc3QBCrhQgK9Y8OvwjeaC0pteQLwO1MFl3z
0ChILp5KmD1diS0v5RigAguHQVoaeqMMmFoW1vqtvax4UECfUchtEmc5gjlWl6iI
SStkLT41U1CxZuTHRuEhv+OMjX7sj6Bz5lipYQKRK1tA2K0ZQXzXYR46cEL06I/G
KVbI3iBeM/Nd96CEXiPqdE6WaICxORbuopZsGGX7SoTaa0aS0Pn1cksvjB/eBSGL
/BCXev0j2+JTeBAQgZ9FVs/LckVaGWugIzlObctSrW+RJwyxbIy5FenAniNw2LKj
xJNOBAw9C/4xslUT5LbWBE9dIfW4PMTVnkI5hxj3PlP7uutyX6Apqailx89mJHrh
bjFTrZWBlu/HEmXpWhaJ+2nd+5ViyJ9Tx9E6BzQ8KK3LGP/t25NZuevHR+hn3krT
WRnpvc1VUZPBknnAlyqgKyIfwgx36tLfN/oY9BFoHA6InvuaxMa72A482MOCbXxX
5zyWhkNKp91+5rt+XBfDsNtDs27GJ5ebaFAFvfIAsE3FmYdgyZq9BK02ScV1FIP7
fygJ4X90WwGy5MW/WyWnfVOD5tjwvxO7GFveNxT6gED6i5cYlf73gdSBJv4WA3v6
92pNTqkhH+4vkjUTX7IIHf7QrjMM6V3BpZmKQPKk4u5CimBgT/bmPJrPzNhEibd5
+ENSHv2XQy0SyJsEIXZVxhhISjbBI8YXlizxXg3hHWEe551lKGDa/wzdpPfol408
PmSryUKcvb6OgQdHqE7JLMztJsbq4PnL/FW+nl2lJX9dIOyRm9GY51p67eRk2KUM
yILgEowiYVCggqawoqFA/6AF3c6juvItZwf5ij8ragJBL9sBbIhtMA2AMxbld+Xn
Azg74McYONQEjcGSeBfWvwwlbsG8JDZ9eZweaJYplhF/31xcPEl67qIw5rVgBRew
e89v5VmWGNcxiJQ1wrjdMOT/Oa0u7X5BpnaQGf89spOz14/P6R54oe3NdNXII8ff
1PC7VVD2dWhbdpk0HbrDd4hdiKeVushlihqA1HIWQO/ORgz3yM/VgUSblpIyT+RJ
C0GfiVGdR/OfYr7ynuayILHECAhJ9ABDJEnF8XegFgMpFTgQ8FNsQ/iD0otn3hKl
FcWqAP19Y+mNVFrkeXzG35qUlf4l2N6Gf9nR6eHxROwTM/wFA+Xq07UyhdSCUtp8
hoR3/BJOi+tNbGzScB8hjjySBQJqgMpR1QvXFHqGaB7ZKn9j3tjNUmftCVHrYCdx
J0iLBKbfaxc7PxQvMFZqEbjFacAfn8nSzPpyvArxurhapOo0610LYw5NA0rGOWNs
8sHjU3GWGHEoFx95s0UwDNkhDozuZLQX2X2o0vm8OVjZMbg1qn2nbFwlxfaPKZjS
SMyWa7XZInzd1flRhDbkUv8oJoiYV4WKwufjUEPdXrVYJe1nJn/ta42xzeF7VsnE
fvi2XauOlBidc7Dv9PQAceahDivGlXxzWekSz7CqZuehdf8QtfvrXdEaAkdhufKU
qJFQVfTmwPBxgzaoID4H6q9GZXkJKuSbAZtUvZkPWkpLJhFrXCB0GUdAYiOG9quN
dXJQIipHA0ebZDNZGlMIL/zFfUd6Tokr56z6mQapVK/youugyhA+zq5g4MiFYxhc
OCnw08FQ8kgR2sGTcMYOtnvzamWamSqpSZ8YiY4+Y93PqOfbtuLIr0Lfqn7UaHNT
46FhdgCB3Bt9IE1de9BFFl8OFykrGFUi+2N9v9B2YoShS7faLf5jXiYnRPDlJaKy
J9RYUlYcq2oazv4yJBXsmDeXuaWSYUdN8xS1uJHWdbt6COg9cLaY3kZPxa4GzQDy
8jW3yF7H1AxoiwmgVPbV17BrKDjJj34yTyeSXQhKDtwDv1BRk3xo2TNyevlXp7/S
iuntjnGo91cE0FJ837FMXfX1kOI67Yh/f+sB0qBPUSzzW6T+4HzG6P1rz6YjWIEV
y1E1hX/VGfN62rolZDOsYUbbTcSSt5TOExGZfOzjh9C5nYrJxRY72UfkyvzXmCXg
7N6SgL6RSTjXagkM2z6vOPT0mltCl7dWSJ9EdcmuzycEPIMtVHc0/udKzqGZwvgJ
FAdPqxuTbgW+th1COqc7yLx8qmOwJHRBwPyrEVlb764VrlfZ9Vu8Q77iVeyTEkTQ
dWmd91+RqARPQb/2oJzQOnXGwnFygI2JW0Hj6KfZim0bsNmIpT2VN1jH7HPn6Lre
IouA49PfKJLjPrAgjTiajG0HJiHo7ymv0huXS1nbi6JW2RTb59Nvxrz1TWku334m
e9BCYAlfcyQL9K1A1+ol3lO6VsHeE3yR2uXYFa9N9F8lspeoyPPUpgEdxJZwrwnb
mGVp7gYvGeJah7Jfy8udS0S/TM/xfFzJk6S0M+O+cvZjaekZwZTiSPmssLBhwwgF
uxMoRpGW/kTreT0nL2D1wn+ZVUZvG0UWfkMd1Jjv1FnxXi+jSUhytVXsegwQ/IHN
Gn2JoqJzNX2LNx9gKqgWxx5ARrM1oOOjec8dfleBd/+3/fvXAlzl/U5CAzfTU6zS
5//vwR/W2E5BDov9AhTz4VIPC3KId4BUfMVUTe1ZvFMHMqrmUcB/rSI7QrZHsrJp
51BuQE2D46W5slRIO+fmgu1JS4KwCBrPuG6/njFIftSdjGSCE/wK9ttE82pvuZui
H606CyTYH2g2U+RDdansjQ+JrT3BH/QkZCsW717qEP4oaQeDF3qkfom/dGP39CBD
JaMwp9GUng8mIA8zoJrh0pLHklvjtys0N6zlSZKkVqdUh9HvEn0AFa2F6/Mzohxr
/7+ZMeXKlmBRBG0hs1BcoIYDowjWgSQX1Z3LZAHzUAPWSXrcTY/OLyPyO9scF4ev
+N8y4q2ajZ1lgD/B7gl1TyGdO/LDSkuiNfm0mLScowYKqmoRAD2HV2B0290Yhgtd
aSMnLg4XtHyyUpQZKTZhivY6kcuHWsdu92O7a8+GZXra8njcuzIAz/C9sT3TvzRM
FfIoAo6aHDXbowVtS0QnoICgzI2o/d43Qtra8o7mOyHZqR+hpJhLmCQ7kLryVchc
CvwXf7En/XAWm9E/WWDcwveo+rAaUkGpBK0JidUsYmMa7apGRohQwdh+SMRwL6yG
d6ZzJap25/9Gf3e6HxaLGxK5QHFzkH1pQdUF4kMlgjpj2TpCedCamPVbEwyman1b
igHXeUiLpYOqdViuVi82SfbFIRcZPlvBsUqd9g93hXy7chvcUW+266woMjTOq/y6
Cd5EUtE8/XEv5k4SyjIfRg==
`protect end_protected