`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 20320 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
YachDS4bpHRDzLXFQC4CtXtH6tDruW4j/a72I0JM1JXCa+dDVGNzYKAVYnnp66G0
jBlqzjOUwPm3jCVCC1xn9tz2ldbD7HRYy4uxPkCHTIo6HKix/8SzUZTdpHlA/oh6
yR811vhHmK85T8Bry2Gygv4Oq9Du8f5uq+5O3Zyi4fVykfa9YQ/IigYNcHRjPc+r
F8SBFwCUFuiJGn8HHsFLt5+NqjHyNn/3QAsqQVTZJZ3BH+j6qTKUFPVMQrdWISbR
VKz2ucW047F2Vpny/Wdd2AKB1ZwTM2vKNms7GvCWdViZDyOQRqIDV5tiFp7wYPkp
/7X2Lk85wkdnA2nYUWZHJqkWi7GbV3jEF7yQn3zAlo98ngbvB9ReSIfd/sIbpv0W
MiSDL9E3XM4hrN3MxZo3VWY5/VfAI0NFoTzdsuDQ34/+uupYaIOigZRbQ8hnqu3V
F8PL0rh3QZWgrQuUSHJacVTvC8LrwFoRyDgVdE0sCn1azYffnc/RR/1PkXKSGLS7
ULj9aI1JSFY37Z57jy7LzAFGR/9twAjrn0oDsoj0DCCEy1xEP04vcVWVLbphZRfB
L8ny5FRN8V4qFXTzmZlJ2WbFPwMXc3BeXQKMws2vl0VBcLtXIUYJCFXUrZCKMQ7K
YskOb2yRAxNZvRH5y20IId6ZHJ1UD9ORC+RoFVSPGJAkOZ5y/S0f4Uccpeu6gtG2
vKyi3umUnjobK4b4rf0oJtjy3lF6oXkvmIj/BCu9TScMkkOyCEXxiPgT5bPXFgv2
No253HXCwR5/d3C0wk4bqj2dIGj2c99eqNHiDl+f0LJW3bdlE/B04uLhuZu8c/yw
02y29MZtd6eodPfezNpLNSKB8RvW5TeFut0y06dMIqe0vpmcPGbEfw9M1XU8BOsy
12AedirqU4SEjF1l4DsAFLbimjRI6aGWYQtGrZ2fMoMGOaPijXVEMt/yGa6cmimV
T0ZEOEmrCCQRMwQ+yox59ghgtyvMaz+LYAc4EanWZ4Iiz5Tyw+r4WW3K9VL9IxgV
mxTle+iek3Fz7aLijvrUeOwdCUJFJVc4I3JbWDwswXHP5kT8mnih5vuowQnOlMI+
vb1csSDKj7PKNnnA8OhF9nluU6dT9UEzHBN8QQjOh0LiRsC/ylVw9ANAWJqV0+4r
8QjqCgvXMtMmqVVBviEFwSFLkxIAa8SfB/6OzO24o7rYFmThdrA7kIZgs6VoackH
AaR/GagcWcqUoh+fBEJH+he9QtgfAzV98vI3iGHyJ5OUD1KU5z1HONbZENqfcwxo
n8GZVbAE0xFghCDKqwWn7QXs4du/022SC7OAUEIFGaAICYUhhBduTf01zg+mbQv6
3OSYWfZGVjWk7JNN9f4wJUOjtBiVv2qIKSciqhk1DenM4kMPLg/YOTLwL7IH5AJU
JL8VtO5owMvGQLqZQ+Tvp5/VM8pRlCHG+8t2tFc7rUf+bItBVmToj8SvskD8tOAC
/NF52qhLPG5Ib39y3OWq7GmVVZ5tcRHvSujehrSwqIHfta3aQzaXkgPczOyONwI5
STELMkMBYq1KDs0TpEsL+ttYcLEL/yVD+a9PeMvWzXsMDjXZklSxGqVC+W8UN0SB
2cLJKcUpjHFFl5FLIRghVz+K+fURA2LccXH5JJUP1CZ2NMron4Tor/j6fKb9a7sN
L+f71grRSK96wFWv6hX806reJbl6wvY54SX/s3ELM2+w4FwfO6t/5viKcEgUDj3p
zxfsNqIgr36+z1kT1lxQjhVMxqNGN5lNj8w6T47L2R1/M0s3EVB9ldRiqu85O06u
tfdzDlA4xpszIPsFjp6AGjME30REMJHK9350qB4dO7si6oA7VLXqL7X1DJgQpFrI
wV9/cczzv+8YaOT3I/pgyolv54P8/0BvEfBSbXM7dB59cqbFvftZC2glQL8GU+M7
+VoYDEh4X6OF99mC8Oaz+Jotr4jOMeRIzc1jU15LIxooNPY7u075BMcPcSW0UKfp
l087wIBGNNu1p0PiQpJQNOwDxcj24iTUaz1hScvWEQHdKoJBAfmFi4SpEwxlnLqP
SXRk6iR1DKz08y6XbCKBunNzpeVsFXXl4HWbr5RXiEHzqkp6Ojw6c86rSALmyEp3
9dw2VUGdW8+UPghUON1tUgzmaoc6hKsTkkUhWwddvmJea+xRyu84poDARY/f22SN
coDTOd7N0VC6NSiPSC1Sr/g0o1kHHy94l3WV87h6TAFH4jcjXQam6U0u/ip9JRH2
dAr7N6G1hazgcaZbrfoCRswGXrgAwVkqrXliTkmddsxCeW8zeo6AahOZXFo0OGnJ
rtLtM4HbVxB5zL0L6XO7JHHfFAM8dklL+MhYWrW7vVqZA6FVtagnmDlenBRurFz8
Gpzg+umFEh3iPCqWn77KOe9qKBL6qVmmYMFvFpuymldXId/fIaAvWBe+aSF3Jg8W
Cd3g7/yri5QZmq91WwoxSiXcDrqAVN5EV0aiaUHqBkOfm6bdKN3DfR4yhQL1MvWD
V+brKXg6B+Po92AIVai2fF6z4xQW030h21EPgXZgZMpbsit7qzem+gQj8dO3h62I
4p171nXgq2PGfZsVr4BkVlDlOZgjEaqwIzni3b9lZnmpthkpzdjTuy13NJ1oFdi9
FJ3hyVx0ZYxz9ik/YJhwhI5S/4Blbgg54l8OiEgRoEGuZHiRaFoHG1eAyrdRPje1
FDYGZy7G8gRDchqEKj4cfmso3P+pfF6GWO+hFhMdLMdtrqweFtDgz2ShjpyHKa1D
R/oe+SgQ2Yxe5tAbWx4gESgTSyx5A/z8BCXMjUMlpdCEFqrqI0LY8cGSk13AE8g+
waJjfPDUYrNMf3QvdDQmCA48ludB+1fY4X2yDtWtUi0t0GvpoGGuuRCOO/fh2y+T
eQDB8w5A3kieKdBxnuLMaTjVt1bJRqLAlgdBdcnHkE3VB5BWZoYGXHT2Kor48/m6
D5gxZAADQ8FF7aUWdrEXYS0VK2g9QO0egECXj1x2ySN8/uJiMb/pezNbtSFbotGh
RU81Jb+MoWo/3uL3GjZZpOLLwitVWsE6bbzKshwPm5zQDo7OIG1sLUxPXGlsudae
v9zS5klVuyQI/x1RJOgxf1jFNm2zF73w131zpHZHfuTpdwF+2buVOsOzy3yHX41C
5fxw149a4LfdgjBwnGEbfE87c5umgtSWlasmEJhgzklGZl3xi44xL8hcAQngcBx4
QgaTcMoBU8stNPqr2FsSTXw3/dSDhugCobndsaaoc7Ov6hMeuOgoEFL2/a8qWsvR
i+/9yYjQIpLAYww3BMHvb7XdfSnJFkzNle9JReMhlDnmPucu+Sgf2zQ95xY69LjM
ghFOo3n1FMAUsOAl3ZmzBoABwzDSLk9I00WbJZlqS+5izyBCsO4s6HEYCC5BUo9K
vcDUcrO7NrBxFl1/jZXfcYFT5Vl4tGYPp4wejZaNvalS7TTMmr+QQA/ITIfYQfec
mSNEUIfwgAaH0foJavMyaG6JgJ37jDtUF181pV0Q7m6tKHR18bSChTu+VniBOnVH
VUYh4V+S0A2ELQRIeka4STEQZ/We6FkuhjJeqGopi6nlTzWHPwbYXJsoAAptHMiC
Z0kWTSj6OMXxcC1IS1uZRGl2M53wPHbfQEGj2pq1ydjMOboEHj/yPcwIj3fNyAeV
H8X7bRkDRvH1dAIp0j7syGF+/DUUzV/d7d39dARChGzI+U8iAN3VUWAIs7czGgES
TKgmPBSmcUBf3EHVBKfVgzy5x7Z4wDM8WlK3YpLuw1N5ruH31Vz8kWWq9ht9u1yf
YdrYry+sybMgHMBvFuWcjJbB7GAABEJ47WWyg3e5jHIt8+LViHEsbyP+d9v7cu97
xozMUNL+ar0dz8F1Trbt1ppcJCfERtK9sPyb+wA0X418dlyYV1ydU20RUmb7pDA3
pbddyIkI+dlETLZlHNRz/LCq51AS/E8dxHV4hfCzZPZSjRtOlfEtoU6xF0GJi4rB
PsOcgQOK2NyuzkfXaFOtz0ZEPijJDIEzzzaJMrmD+3IgPmjkBfPC96XvLr6Sroax
hX28lRSl8VGAQfS6sZJ70DN6Vj7JFE7o/CQdZMJBHkXwfGI+UKDsve//oLHShjxK
9cWE2CFRcdDgvkC9bR4MtivcFyccx86xA8GykmLQNfZR6383/yU1R0Vw5GruNBJX
CeUJy7Pb2R9nlhc0g+NhCO6/OzmBEbAy5Xnqe5+hnYHpQuCuNh7StfPV9dhe2FJ1
9PVQOd8sMUjfW01i0fTK+zEP9ekUA0euIBmPSnJWMo3v5sHJryrDmOsEdxQ6q3Ql
3uIMP0CRI7Phn0HkB5IoRkKQT/ijdkzg94MmyEAMltZe4StuV6JDIglhauvtrkcv
ZyXzjskGWK16OM+FNKxhYwSYY+RrrPKg25Q1l0C+P82h0UzZWntDhcG0Rilr+agm
B3zwZhhdVahMRSMFCkXttgYm5bfpLdqO7fgut/ubjjxsfhWxBRkb7DLdPxNHlOXn
AgA678DCP6A3Qrp9tgTfSqbUnPfCiLGZXWol7qZ1/UTmCNS/u+A4qmzp+25iiOJd
eTk9+wxGj8XeDXR0+MZ4Gksn25UvsbQEGQcCHWMlmvWjGGp7OEztDDez38jRgSDZ
aK4FfAPgYts5vDZ8WCbkJaMHiqVkmtVfrc6rpXxvc2tdYvavGDIVSN6bIK06pPf9
7EQG4YJWi64QJAnHhDtFkC/CvL/9ENiNZp/U4S2e2Nneg5ynv4o973uZQCYRbv/C
KQxk8JF7Ba/EzsOs3MsQOaHXigNGYQs6pQU0bkhvYCHnQV8FyC0eoro6Ets9Fu1O
T7mFwo2/TpIA4I81xJCzxvK6VWROUpRqWy+0EIAiCYMpPaIt4k/GX+hlyYAEvCBD
BjiiCOWAiN7HcZOebm/VlyymkLf9bMMs6CVEiXtfvG0BhDcKhGwKyL1Csk+pFnTU
zvUNXRbDcVQAY9eym2eVKINZPhoyWAH3Whp1/2chzhULMGQctsJG0ZHRm9g0QE4v
gDLowtYm1CL/ugxH1DplYqgCDweNj6VpkY3T4IX/YWlGu3+iE5aXwskoVo5YEfK/
g/gRgMTaPgcj++gIuktLbMMqlvUkzWxIrMdcT99C4EdGtrSS9O+g5CxOah8AhwtL
ocFAxFBtxXvhrycckxw3CQqxWyymyxA3bZlTTPrFakd/ANaOqAzLrUTsyzPc4P8v
q6S2OZav2BOkj6LFKBi39Y70/fdji+VSjeAdDhPUO9hHxj1Z7eL6FLY+yK0K16hS
JmZFOajA8ozyb5m7EEtTNtoSsFoC3lTa2/GeEElqq7RdoSStPTYFdlmMtV26850k
YJfJOgG7eQb2xUVKVi620ANDyskgTtD3SIcNoJCelcNJkWPjjAOBI4dysAMgy/c4
VjhjEzobjkylPM3RqAk6tc03EEvY580r9Bsi/mjGaILs7MIt8o6ScBEikLPSZBM1
XhbMN9PKMOyi7sSgD1xvXnGDXgTDjs2/hRiXW3HXfzfl4EnNwkoJzwji7E9znIiM
eH35glDQrQk1NjXGvnVMs+uCd+hw//poscTr+NKHyDAfIdV353HvGAKa8zcg5I+C
tWXpKfrwpkOWKwOE9ZKEF8Zg5JLtQWrwSGqsGd5tCpwT55yEXP91Yy2Iqfw4Q3az
eNkU0RRukbdRYafECmkrkW56creqhkTY3KCSrSCDmVxJAxxx+VStrICcaHWKcXmx
f7ChjNKCTBZeBrrCx5eRcaJ64Fh8nc0eg8vLmNgaPpc0SihZZ1rhB+l0ZnEzBZ/P
N2xD2qWILst/4A7S98NtYER0NT+X95pouwui/x8mDOFwD1OLtH3eJ61wg/cUFzKk
OGnXEa9NJa0tuWseWx8ErtHVpRbnvS23J3rHGkU7UfrAA3vZNl97P54jc6liILHa
t9zW18exSdClL4Ju1lRdQOvztR4/JbJCdh9auDB012Zstl37qwpBL4BdjRK/htGQ
NSckGHkn5uKoiakxkBzHIckmArrL4FPoiee3+MoGiCYi6Od3CsoOl4qubQReoXT7
njeq8QRw7NJf/1gRPusTEck81hu4Ha9K7KHRsqWN/Ffw2EhKLyEu/yjNguAL+lDl
un0jq7nopB54gZuWTM/9D4+k2PHY8uGJkmgWBkbpkpGTAO4dSDgdRAqwjNSopjES
tf0reKv7ZS6Ievj6qir3s2PnXHut0yVgIIUbcAXUN7AoUWve+gM+cB8R94b1/2Up
Oyn4CWUe+/cWizG6D49VKgUINFtewmoJ0JThm6fHJSbiehEe4hiUFDPCR27UNV/3
KuGFHjCqTuxDERf9XH8VXv/dATRNXCpAtnmSxmq3k2ORYAx+OndZy8QRfS2qkOz/
gZjaxqezRUjUvA+e5IspiUOuJP3/ko+qe2Jg5KT84ghL091ZyZW2mzD8+GDFqB6T
oSd9AFXGfNYjGepfopLNKMufYH6mCGpLsY/Yoi+VaFtQ3tKbaij+pRs5mtlrLZxq
z7YkGJKk2Lhf/DwWRjBmPi7Vf85HVli/wOrARyP2/3DVnXRJfzvfSejIcTbo5XBL
A2ncSPENSyOANo4FhvcfYUYRSuoJC5kZmri+pP2SpGm8O2+N40ahYydfsb1Fvzm0
LxjLhIi7XLbkapRkz0fT6zbzqrAWXiCDh3IH1kUjPAxbh/gsnldVzLweBpsbXOrY
HvAzvvRzS9+BbyPQgyoltiqGdJJtc8hPQ0SVTo2knQxYt6qj97xKoeufeP8RozW3
FMrEaY84oAtJTiJHrnGwHQdkjh/hFMP1pCoPMIKV0UwPcanpVWkGgjJcyciHXkbh
YM/Jzk89vSGqpg9DQe3clA2EVXAOw+JQUPPpimhKB5z49SVh45Gx/Kv9G8hMnZ3X
BuCvd5DFaLRoY13gml80xPR3S7LF77TrwfZNcNXRdfjSgehUYZyAog3gfL+paIPK
iTsujy7PzM9yDfW2O1EagtqqBoHoMWP3o93NfIGs7wQGEC3dFnDuGRHBc2RAdMPq
K+2QEcnl8SWAfWF1UqCECiTIv3d4ShptemyS43aj8yfaKkqdYyoP9YIRpxyIfh5h
N2qepeqvxqad+aV5U5tQz4obKjP4wUus4yHENWfQ+HVkqFjzpof19I2WsTsAFH6M
mToWZbclD8zlB89oknVzw+9HK1j7o9Y2YrT2/IUm4EG8zf+EmWQQo/56sKJmS912
j2ANAMjrry/iHzjp7NqVLVHD/A3m47oajIgi2PEd9A2dEXoEEzdNEEbJwC4A+QUr
SxUwBBGRDJw3vdDcrd4BoP1vvKWsLF+GU9ygo38iPEYwtuLAlSXMlomEPxupGduD
cZ/gZTca81meC/EnUm/mozm44f6C49f45DGtr/zyDX6MMDgQ1XqP0hFyIWdHTfCe
H/5OeuXJYO3XSgkkchSi8yXPvgobLG0HBQy1Zu678aqu+qimQL1MwXpUFx9K2JJ+
Ft364fKjMt19362BWTfp6kWw03L2u+PZnpW+W0Sgwx3dBq4DQVMTrZKhYCrQnvNf
iSNyv7+SH7IjviGkXDbH/5ROvWkAIZyjLyhJyYLt9184ddMimfKv9TTChVUiFWq3
8BbgYryZezkuMA/Attav8DitxEGc6xwIaR56P8+03goZ/6WGrFR4RHGBVlZYzfGM
8Qul6DYF5uCB0QZZo3EZJbMwtEAP+BNIoh4vnR1xWVeSEM6SPEuraF4TZ/utvP8l
+wu2T/4vJC5x+Cv5ZwV8ARgQdXKDQj1Fij3+akflTOpHnLs1iOhRMhXQXEzhMjf5
Pa2EhgnsdghNyIYuMlbc9H93Se27LKCICR+ivLZpm7T3HZeyfYpNlGiYRX0sGnFr
IE+XF/EMzBr93KYS0H/p3401omR6VY7H28q/Xpmp2dFUWcU1WQ0c2Klb0r6jkqVF
iBmKLsncuj1fC+AWT1rCQEpqxBF+B6zlNaM46KsCBci2M/+bra1gCC56xSiJXQmg
deOdMxLPmN44oLGFhtBucJaY9N8qFSAoXtL04QasJ3bOMROlyJ0CBmujkCyuGpap
WFLNKepOTjJ6hqsflL+uRTn1+dLmsgD8wWwHdqi6VttmlTnico/eGD17L3kURu+u
59BMllkZhSxw/nqa4Ab9Xuj+GrzFPb7uSQ6g55VWWFz19smRRQDgGM2Cf5FTwY8V
Yz7XhWT6PQx7nDXae2po+G/SCRaaQQPG5RKlObqrucGOpL9+KTitsw5HHB+zlBi+
tD1GsEgZA0WGwIhJah+yGYC3Kar9nbw7T9jn7wdjhDf0Gd6fU40pTh6tjVEe7mZg
XAU3eLuSGO/Of8PkaxvzZ/upuBsAXIXfI6h/DrvsVKmUnw4DlWQ/fQ/22NTngF17
bl/Vu0nZoiE7KHFnp1+6WwXkg3Mr77UCmNTmXP5c2bmlscSDpUieY/MFs6IYLC2Y
6Boa+FL6rG/0VaH34W9+lC0nUlYpV62UvzHa7o/tqo/WJ1g3/U6/cCrjSiL+Mk9s
znZ5PySIwnkSR7eQrawaX8dz5s0HyB8N2efBdoN/GOH6k3XJ7uolqla2g8QOZlZM
uXIpEBYMUsmKYNAaTxZnR0Fe2GqW/yhNxlmtQYRDN22eidWS4QCu9aeKg76vCsa3
0xIPHy9XgvPK0SZonMauQlLiV3Qnlth6xW89/dhOlycvpg8+zmLC0/61Kg0pTqlG
6eF0kDaJ4+OW/ipJF7uOZfU7l6KhlDOlZJGpnKBMvuV10U+M5VXyghbplQxcNOJe
zik/5RvWZjxF/GlzN7x9XQI3N0VU/x4DsgU/KysdAa/TrJLV5pdyaXquOVtoz+t1
Uxqav/mW6eLe6d/x1oTXywC5wCnkrqkfkWwFnAVyVEisNL8YbiDqunVIzSamHgE2
4/brGxu7Ks0GdOxh3wBbsP2ZOyGfWlUs9kZap5sWSFitJE8Vbd7HGDX0HiSettGG
poo2WwBTMnjUT/Nk3/+nb6vbqoQmjCmmaPH3ce6l+doT4qAP+tn9cSsw+V7oLAou
An2Rvf5zJoEq451uh082O53g8btkBTNl3bcMqFcsAnOCsuCGWi2z1VQIvO7M1oBv
s91DnCmmsH4FLyPkL1FsLpsFdAcVkOgfHxkMUZ1vbmmULkXKQXRRbG0PUMwCYV9G
zSiRr7HYM0ANSrKgg4G7AHuVG6sqguobegPhvcNPwKLoY4m/HRL0YVmeiYqX0kUA
H7R91rpbewWNMBWMwlYDw2pkK9dQWtC2iK7vGaOCZeG5aLQUI4c/+jiJ8yf6QdJd
Iza/kr1l+MKzZYfFhl8kQFPd3gPC8/WM1HhmgxnfnrI3egs9dTDYCTmXXGoCKqFG
ndfg473LjtmgB3nsOGCfs05cBftfQTGxg2No+LrbWrdMXB8oc5tsP/R8YP8v69jp
wgttzF9Z+PWvKOHXk32IL6ZPfmI4aKN3Bnw6uE9mxFvkHW+GFCgJjgZI3vN6CtV/
gJGBblrGr+IwE9gLL8rqT/Q6sdmixKTeCCRP495VWVoOA+HqPm5Eb30tSv4/G+8o
LtWlllj3TQRFOBqOHU1xu1xqw7I6ciiJck3KMmzxk52QM82EdRtw0DQF6Z5gqwR+
9Fq/OnvFKO415+fpaz+OZ/177I2nx9I2+SvSRyPEU6YD17rc9JqOlCQCa5g5COl+
kFjWdppHvLIs5fIpUhkKoFmORWE5nAFB/ghK2Oqk+3S4zYI5WdZUqlUZYx3pXHvb
0qxGdBp4gTt1CZcsNUuOwu+vhROVKROjJcbGBYZTuaQDNXQr9QNjMmeGYLJb0hXT
a/0vxw128cl++i4sZxNjYc7U71QlqzdB9X/WCfkUo+lNauFuEonBqKAx+Cq30Onv
0e4tEPQ0QEMFZYWWyDx37XmHMd5P/WDFmLEL3ePFxkBb8KX3HQk+HcrHdwGXOfTa
g78HtM+UK6D0bdLb7mzEsha7Aki8wS84u1dwLhp8QYB0ws6M2s1QBsEIwV6jKy+I
ftPEyaI2eoumu3A51qfHSNT3XU9Q+iV3Brb7cA+ibLFxeQwEBUxH3gdd2rECYX1s
FVwRixtivFUB1EkG21DKhnZdWGeHUaCCv6jwLfD/G6eGom69f25gNmBKFiFU35d3
VOiWQrHKJ2zfDlAgVNS1HPaDY4Ezy+tIPRbkg05aw0RuzLdnFulcb7pI2EPKTyYB
XscXIm8Na5M/hu7e4YD5IWv+hvgKKUk13RS74USgmIiEFEbZJGKSO0b8YGOXMdY5
JGsNy3RQO4w8Uc42yJrI+c+/OpVxVzTLd8ierwPJgi0Dz+MNZICG4y8qsyI/lB8C
Bm9o5anYga+RPgKSxTpXfneQSvuM0m3v4ToWVtRyFhNKk8tepL+JKNiKAiEOTCci
WnvdYsG2ik5WLvDVxn/+O0VPzaVB5Tgi5gZw1mhUFcGp6hCfATnb4mg3qsn11Krq
VsjrOPrG1LxLiX05QNfpQQ2R/lv+fwOaz7xbqGudluZm3EHjRhFCo4peTwWqme1Q
BSY9A1tVXzIX8oisDghPkjo/5eg4M7A2qhLy8aFM0TYDBysTSN4wsUdE299vbcOb
7aUZja5VXWKSVoNHj1JXj8FjCP6UJGFP0DYtBm+rI1+daFuMf6N2ZOCiL8Fre7s4
1eSiXTtF9UOR38JSHQPeP7ZQG+MwGM7Uc8Wp5lINreL4v1rRlecbgWQj+ZLaNcuL
XwFwYPZso6jslUJAE4EHLV7eiNDCZhRc9b5HixAWNzBb7u2KSq8viDYTA98gd2HY
wL2g+BxHPZY6tnc7pCklIXJ8vjKgowMzV/TSqMJ9iE7SofGtAzNPMqpKLl015NIQ
lTsSYeg2DnGgBrMmdZy+LonRoZfAnElrco2k157j2qDIMFeHifENxNIgbv1Q6Ha9
ajx2fxwiDhl3Jz1gxEMG/RD7xgCp9lq8y1Spy9VAxwpk3ZwOaRL8kyj3JQLJVdiq
0nMAP3GlchXl37Fct1TrTZ4oBDWzd1c/tOa4D2kEynMwOmJ8VG5GkFaHoovsmEgm
WOJhuVoIQF/ZgdJIuPvuFlu5are6A1sT3pzhUNP9EKAAvVezSnhj04ho5IQQdjOZ
nIebfR0GQMroenClEdwBdAWHPSCPv8ZGike6BlYSgYKI7YcaZcRbv077ya+PMxf1
bFYYrk1XTfgXjTs7VNDr/KvzTJeu9QjTS8tRdO6Dlu+EceRtZq9LJLIOjjr0MwCr
qiMlRKSLfscvy9tBTT3BbBZ1CWr3u2l4KgKrv9gmIvTb4mEcS28DE9Y3vL0Yzpgy
LEpS7qQt95EmUgHjL6PjyYrHpmgwLRso/3o7A14ek5vTXspb0pmu6tgxM/542+e/
+IxywbdJqlFshsT8Kl7t6Nu73flgzGC/GSWLqWy53RCyjBI3LQ075901KnyuEq8D
8gjoa61NfHUlrC4Ap2ijPQv55QPfsbPxdhHBIN7YVMrNHVhDAKVrRMGMWJIlOSti
KjaFLiJBiRs80b9B5C5WoAerIEThk/A7sqcY2uqJTRZOJr/daTQonIvnvNNMDcur
vt443dBguqFp99IeurxywV+tN+XyINRUZu/wMgDpBFABpbrwF8lbaabsiAdQVmb/
hJHftnybXXcPElZb30zQsoV0KVsLJRSVLnC2GDXUywHBBZU78M8aw8vofQXaVGu/
cptDX3rtSHFZqn/YB1B6Ack3qyy9hDFj3JdoviwiAs1yY/IJtSdaijOuww13/U7k
yOsju7W8aiw3BtQ1wicOHLQrP+NfNMUtc3F4hEe/fKa+MDIqYPdjAlbJR1LoyNYe
Qn9diTne4EzG84YDU+AxgA9raWwZTOYT5DFbiFR2LdN8OFLNJooS9i+tcf3vr/Da
Fu1YDCCA5vGHfcDcbDK1ylJkWVPvsfxSZeYAL0DW0lzoTYtV6JpJz238hPS/pGLp
pQw83gGFE0JE3fAKBsFzgUkPj8rq2b51tFth6BkUGhIqBGaj+NJ/HfQYGjATM/8e
iZMi1Kp0RBIaqmepwaALmOhTpCCyA+icCYibL/9WCEaVKZghws77sumajnaFc+mC
jiJnzXxX7QJRJ7wJ5Ymjx1Fs7dboI55h0v118PDhtlHyKj4+jUiyQLboD734/t2l
jyYRGDE6XytSPbrOd+cbebUZOzHywV4YUj4PIf6dMadaf01J+K0Pnh5bGyZw80y2
yUT2CWj+7sxgQAxg0XQJx6goCICM9HIw5Ei/o6XoDCoaZnj3rgEQvI41lfhQTc/9
VkPUxxiYUwDcBrhYAho/AZoVmcEo6ivWvAqMBZspXJ/w84/Vc02X4DH2+VbSNEfy
L+t448R/OuihFcRHssH8ZQ5x2Fv+p3bK9L3BGsPcmycgWwUcEWsF9q7UVopDGMHH
hX06ewrlowgmAxeTvlpigx1H1szt2YX+mzEcq3F1lbGvcZIrXDzqSmnb3QRhKXMc
U64u6PQsvu2ho2BzQgv/mwgl/X/PdDWXoAlHznC1kyxo4BSZVTpvNm15uuPTGJYW
peZY7Lyp53O7M8CgozQaGytA09pySNZ19G6DuQ3g0sz0LdRlTps11n3N4aTFPSNu
PlmPpx+2KTIXhC9SgIVYpgSv5VgOjGMjxeMdFrxiq6kZvu2ouQACkpG3wyy9IZsU
Ks9yH61lsWz7PEjRbveNym1rYySFlYGBcxmbZTXchyxrKfHPQd8sY5RYXr3aTpQH
/ZY63TaxISVC4rScEJO21oQaJg/tc3FvnB9MCdjYcjb1Y0dFf+2EzlL0MiayTrY9
Pd0EWlsfj1izqjAtBSBvqicmmS3HhzzrtIpL5mCNlsNsd63H/fXQFDsFFill6V1+
98wbdpeuaGYTVK6xXYdFxsuws8cddc8MH7kEI3oJ8MNbr6bpczcmZS5vbK4m7XyP
6zQUypRdpk0i3JftKxSF/6HDHiEFMFhtQiYjQ5Xev3rdSxPqEiagJLUjKwY4k2xn
l38rBaS//47icvtZDsSWQsvgLF5P/YJpp+akemuRy6nkNVT1MuaT2c7HN5TGGGC3
8vhwwypOe7RsnuQ+0+e1lYD8Y8HxFwxUh2jlqHPJ07ewYpb056wNDSKEe9uEmxYN
WR99NtGzWcdMitGPEp2e0j86ERcarZiZa2Tk6LZ+75sJJ5Zy07vZmrSEZR0pEH/v
c9c3aVsR4H+NOkE5aiWm0ovfV9WqnhH7BO+B5a6HkquIYbrjHtHFRH+jQBDqHY5k
BIJ0QwufSn5PG0s5QRbU9Fhtj+xGc5faH9wCg08w4qnIEgG9VfZkvX+JavKTLKHw
l2moBHkVpiF2cO9H51lMXuU8hOuSQxv7RvIITAmagYi5qBsEnAQRk3SFDdZTVPzs
ZHT0fCeIjH1jbwozmWOel49IgRGMHSgnpePzvkFxV0Z8NG6HGWmV1SGU+7PC9OS7
noB2FYx1UmSgbFAEETdFTGKHHp7NKc41bHwKyCNmjl4s+MEjcRjuukpdh0CULjvr
zPFWAJ4vjuvdzYbla1wKQQvJkXoyhW+qKcmxAETPZmGTF0GvFXKSGLFRX4UInWkz
cf5LThb0mInuylGaNffRgUgHpvPLfK0s+K8NAWyDr6jo2+duC7xToXj+tWbns2qq
uORrYM74woi+i3PZ/HE59FdfXyV52nbqj5pKZdtxdikwdZkcerrgJ8cyW5qqTWkr
ic9JEtKLLjyt+I92whl0ZZIwORaY62kw5AVN2W0AO4kJc4pT43ScVwUEbzqTE+Ha
+nRIyspNsqd+6yzrDD3De1F5kROCAFbGrMEIUK5yqiOeeTd3q3OH3LS9kpjjkC2O
vqS2FZCa6Nqsr/zD3I1GsUzE3Ty7Tx5qO8qf1kWr74mFcOvrN1xtNN0M9Olbi+bk
WwcbXTvok2oEhsm7smqT+NE2XdhAQfEmfvH2L5wSajd/WDuOJ4pb/0oTBVDj29Un
VmGFR/vyFad0afH4uvR1T5ozCPiRGOTdWPiuXZ01iokP7RTQXSAIkKAgKooA4ouX
1E6ZfroX6k1AmqA8I3YLId+pumXyiRf5qZYxNiFuYZYXB2BXG7PayZZHKkn6KIp4
+DGRC8XWawZpt0kgMRSwWITIJo5OaaLhCIZN1jSNUAMJlXhnxNSdA1GvXAD41fHp
sF7zhXxe3s1K0Bn/rk9Itxndpyb8tQWKRb+0bOJbuuwoR+XfJ+b8xhC/oG4/15PO
las3WIiuIxjBfZwM8U7kBcWis48JA/PZcH6G8EPuRJiV5GJNi0kEpT6SuCVukaD2
CSkDfSgvF/8kLgkRmgz6lXG2LYKN0zzZo/gBN1fBcxx069quESHPl8sOQngDgf9x
ucRO14zHABzGUsQ4pxO0jimLSJYIVWCRRcGdH6O6yRbTU+YZYe6coLdGnbFg5jd3
ppIlFDuuv8AT3qg9e8Hp5Mm6PyvJnsGGWNO7mvoadNFB2nuBYMExPLSXUe4n4M+b
95KWp/y9N4/BtWOQwa791tvm08X3EZCBOriieYlYawfUzSLwpGJMlGN0MJYcqZM5
tlo78ZlNicpmohVfhJ4WY/MLR7RU0cnlDC0xRJpSvG0h40PlXjHj/Uqu84rnE49x
OG7w9xSvY74nTNdMh2hzPHNOJZdQWI1pwD0LjnYUkBXjkeU3zTNy2qXbngI1G1Wj
Fek0gB+XBWE3Qhkz4MgReJfItA+TR2A7Kar+BxQG2CD3OQlyyp+5VQ1CV8bXOrbX
XccRit40APwhPzFIhi4l13fZfwIZUXkVlV4LVPFLkGHIHXPcFDRoZlWdZvUMDh6T
WpB/tNwIjLlP5FFpQZyuDPbywJCGB0E8MBcPUjXcGBGzEyc+fewB12Aq40ExNjei
pY8vfuTqM/0dFJiC1y+HxQo4eDidpW7vQf9gxMl4GQaNoRVUtgipycFPsRKP18j4
EJGzKIMzXxzu0fEipM0owbtDBK3RjuKc2LK7q5G70e4cnpdC4U10Q2EMwogeQfxg
+DiV84xSyMxxdRa5ecH1bYHxVCYmJRbPr7B4MOYSAtve0SqgkAV1nwA/XAyTFrZ/
MQFkcQ9rE5fDGI3WqXBRTNt4nfuaHpG2r565eU+IhgrbtlMuX4RNjV7qbYZ0au6h
KnoxnbblrU4Z5MDQzVQRJSOY31pHON419ByqN5JDTmVwtZwblPp7o5Kd+KsyJj6U
mhG2GgPIdhfPdWVpvOecv2LqGKenOnSscTcs2e5QCKFVfmtRXugeNXd/JRQRbaNq
mQ/Wsw4jFUptolCEVnQa68ZIf7xO7JGBbd/1nJNdmSQQyUDECRVAzdb9af1DCl+N
a7J0ZQ49kEYsmHCe5e+M52Lg2O9ET98qAyFBpq3i8a/vP4LHlhQMuYdbL9JGRWOB
xycCUATAkzDAGwGgoz+mNA2BP3JatX7Vq9vxMzl86PvUM0AN9AuU9U/JD45v6pUU
1G3i5dZ8JndmfNqX7j07zNZ5/WxxcbBMeJEkHIoZhYKEoZeKb+4PK6mU3lPyVz8i
iFmjKfLa2Wh6TMPbqvKFm6Y4y4zpgJ1mARrUQ3lRQFbx7ko4o8stjeJ0fNb9Z/5L
6DPh486GbXuGw7WKcEpvpCeDOvENAGK6/vMSRIaIeY+fmCot7hQfsN1g6L44ncvo
t2tpKgdOVJWfeONBIgDDrqBXl0T1qZK1pKSArxfkGPHV7AOPiL0GPW128Lbhx5RM
jZFy9cUX3qzjHB1hOOnoXXRHxevl2n9KxkQljtsimkHT1u2L/34/B4Cg/+jVQYYT
Hz9sSeCu2iEDRBvdXIQCvBXfjjFq13I/II1ARm+s5cCYuM7TpTa3oCaXS4QeEwdH
vfCHVZirijhR17HYGIbtIo7XLvZzQFzzMOxeSpsOb27p8pGpKmfTc/kYQqpiFAhQ
tnCb0q/ERZ393u+uaqOtsQh0Ey3Nb7DjBJR6eMHhiwGzhliQdNDVfMVdzPRtwEXC
I2JbezOYoy8ZHindfytxSh5zVhiPBqfMOQoM/IYX37scHBfz85+ZW0xWpTDrMiOB
Kpml/F5Eo41Obzys4i2OlST2fzsSkBeFAGbozSMcQ3adMAXRncq/H6gai5fjMiVq
QSNCjMdkFYTP1PWVT0EfLFMWkZpEGSIfbWqOOD/HUS1zO2UG1injQ+q7FA/vMjFs
MPkxzrCOEWfLHftOnASCc7DcVTVs3g+xRe2dCxvZQVMi4+aNdJmlUYxMjJjkiXqf
mKpmRk7N5GFeFW7hGsH0QwKyWmEWUlQYh5atfkmH5zZgu49L38FaANXuUrnfFB8x
wA2TwUtXkgk13jdaNuW4yolewnxqoICK9rZaDOZyJ7tLvBfoIxIAw7NvgYNTMuBn
H1j6pwBpsoN2L0t2RlOrVNYflJw7Gzih9d9oe6XHsQVzJ/FBCUQv1JhWh0PtgwAx
uvxOtx7Qc9OtL7uZo3cpE3KSPauigQR9tN8wA32UxPMQZ1g1zPuYlY4b2MBdr+8i
FEHt5Y6XN3VZLSmIM2RxqpJn8G94a2KHiIvaBL3bVa3YyrZRZ2HVMTfsNWucYDT4
CD1VESr+32bcOr/2zDyWMiMgfkXIBj4rmvFs01ZRLRVORRK3D7VP6Um1LGpy3tps
LT8WuMxbPbu1MGU7A/jDazhUArEJzLNXrlM8HAkVCdBwlt6n5kdKikMzMRlokDMM
/2hG4NtWJ+4uaVs4pt18YsN8sqN6K4q0Pn/rEZ81/2nQ1RPboMTvl6/AfeXelrbg
90noOMgHF+XOJoRWtJARw+LrZx3BL8ZNcXMt2qaHV0m7jhk+cUNYyW231BWQoj0D
hiMrZb9nd/buFJtQr/R5XMRr2FRED+JJt40y6XO6CM/GffSxquupkNBllfKIqhun
jX+mzTh1UYIJOM58kZE6bwC9EDVSYX4VROju87w5szngOzBmOnFQRSRdG51jFJek
AZu8jXgA6NYAX+IR4v+erw7SrQBLcMvopbCIbpK3Tqcp5OwBmTnmq+nj2NHthsmB
8SgRdUHblhXgzNSmRFXXuytLfO1c5xjH+vw12wd1mp/JG1pBw0x9TvctAX4/ztp7
bjVSlNKvt0AERFiipRjcvhoQ49vaarJJ2hhMZz1zSlSi8q/qXYvnfxd3DSv2NlWU
SYW2hIvJSioldSHLH7Qu42Xl+YnrUfInWF8AsVQYJC8KXDj+vrXEZ8ci91CV17di
0mpG3Lrz5bhY3PaNMRIs+73F0qISkgItgFwmhkrX827KDI8ZV2Gd0I4gDUwn8AFN
sb0YDZhStLVrO6We1dudDYdtMgcOg8iGqVtfRKcAugXTd7JpA/6JFLkKMgc1k3mC
ERLKJ0pBo9rmCz2wrcOi/FGkfR47Tua31Z1vhrCARQ/HRtSKbHdkdAWmwQ1pUZZz
g3QkSHWLJoBQJvUmbdBYQP/HIWn/CHfAS397OvTxOTP4dOErHHYuPPq/ES2Ihvap
mbJCNeqkWza8OY1Aio0NgqHHmwSuV2vyizpq+3C2irr6q45my8mB3xwOxe2iTb/v
2w/VDh1NUWEgDaeirbCGG4EKMcktW7UMHrkvKxdm7cxlva3yZ/RJ88hKsaplF6es
C15zP4N8Gp7zKizCEkzWRM05BK2xbLM4xyFWf+q0oTjLv/3lo4sQu7s43QqdEW9x
2UaUvDJnrwdWMBiOYvWGo7vZYiFYOsI5xXfy/Auswg8Lpw7oUHzuinosvhOByZMy
sjdzXAXwAlqpfRgtkbf+Yc1djxM9yHMeqnpaWgXTSjrjMTEZ59YP5fJ58Pvd77Ea
JNBj9ltp9p+qHuXm8bhnN21YXSWqkVwi4Zrd8AgoM9piZjiBy7K3Gk+zGeXV6/30
iMp26SU5mfYfY/S2pkuvon25TiSVbExhnZ5TfkShJgQd+WR55gotIWM/jNUyUK8z
7+eA15KXHdoocEjP3LjmsuBqpDO1Ppfq35fbhFA2pe9bKD8/yVDIL/LQnqacxoQ2
gxE4Ex+bkPXSW4G/S61dXCRFnA7GnFse3deSWmkIm5vnsv7G+Dz/ZsgZeWZc/Gxg
EkguYm/tE8JyF4jIPRib/73Ob5mOleE+5uPB7hThPUUcDNEvRLkvogOWvHpx3l24
UcxlGFmJe4p3NBq83ItrbwjJ3ov9uSscDnVUbXlrLIWBx47x3uuZhlkEIIwh6WOd
w9ubYENxCCY5evCAr0z+GjYZIWVtMRJDz8q/OJ0hNg9JhZR/LtLg6OnJOTDXmCI6
u7/WVXns8inM9sbrSifJyE/fX4HmT+efgzSxHkRX+9uYhgKbDI7IySLsBeBEi4vQ
ME2m2VpsLNBRHCxbvgiCUj/G/CylwK3LNFNy5IYGpkAs6F4/aLBqINnJU+Vuscz5
4uwKKXrhEbkHCRm6WWSQTbO8cySZfK7/TJlcsInRPH9nqQ9b90YnFDl7331lf9kP
AE8CMsNrwXpZMzGiL7OQ5J1j+8ADfyROjpZrUZmYoc1BfRHwmY6Qqb/OJFLOElOy
jmzK+yjzQM3NajdP0yn4DnByTr0bEjtD2k3yNhdh+Vk1Aa7yWfElRrcM3C7VlNtM
jYhsH/9jGG1Lkei6IIAVc3rJ3EcQWdm1RaV8qJdfn5oLgU0+GW59T4AI/FAq+/2N
ektr6vqBmg3Joh0wpN9Ja9pmYpEMhPR/1aXBDvf3/jivq1nDWkqoNSfZMfoDhKjs
QJVYPlQuckEJBG4YxvMemo1ysCN4wyVyxETT9eVU74O2zh11nawdfH6WggcDA0in
n0L+V83alqYRRP48L6BBRnNqbWkA41iU9nWeV+kbnVk9v7v+DrfzGExHxZlEcNQh
XzpHXUtIWiCo4O9/FvTS5UywODpoawG6U2dhaLd61KsRMa5f4bsiDH3+/VOJsoZp
0Ui+dB4Q/QsMJrLybwdUMrebkDdLSyvEoSmRkZw21boIgdezWH0L5FFEXGh0FYWB
b1+dEH9zjzxOmbdxa65bWcmrA9+mMLs0IvHyLR6a1QPX26bapGSMZyZcpTZqe9OB
MNG0mU1hNwEy1ZiskZYEra3VVe1ZYF+VnmtPV59C+P1OHSaiKPh4X7WO/NAruD+0
dCdwa7DUKguGuEOPpgwv7mM7DIbhOap4TglnKL6oVOqrf0heGPjSX0PWUAJZELx1
20DpQUaNY7aHCFkhxFQ/DNP98EXEwt8uz8K71VRK41lrZreE5vCZqAwyEWypHPjr
u7VH+SgTGXo5pzJKMBwqZNa5PnAesti1zCZrQLYJbTYWv+6x6lmQ388ewcIBZhpP
2iMzSdndHmnQqoCV/JN8tMU7CuIsVK2kgjuMu9dtDnWNP/b/zzGppcOWGTfX877/
lxWG2/TofHN7UoivH2fEuJtzaWBtjTk1+MhBWLG3l9xl+mCk70n8k06HXbiiTZzO
liVsDZ8XGhDZcJFMPH+LEiuQCDIZDGUOM4pfv2MnyiRQSvp6LRxiKwzf+Gg/3Rwb
oNpPe/L5E5laktJ08ZwWLhvtKmsRGnYt/pUl3/y7ceS956Es/4Nw9FDmUYApj/6m
9Me09HbtNs+mCSb1u9UYlRGQriVzPjDw3PaIZTVX9Tlcbs9WoyvtANk0LqmSrpXP
CJ6qHuBeYHMcH8/oe2t6CSiiic0xmFXCqBYuoz5EHdGNYwOCFqx2dolcVR8V0PT+
g5plAnREw0f/pB2pGOAYFcI0iqvOv1ezgP9eGL8gPAp2Akcjo72zKNoImsOUAxi2
1dtfU8jZeofwBQuPyFWjRhITRtDxd5ixkMJFEg8Sml/WzMjLV361D0g8egTRKWPZ
dscAZFQFWKwemZVVpZdkbmlMuktboVGZEcLmjqaCgq5pN2Qkdw6+e+VamkVHiWjT
JIDK8gwA+7KJH2Bqh659hUsVD+tY1rCTsAeVrfvBKS8Qoz0KuO1hWKvpgW41jFvu
9ls1vmdLzzVK+d0P3es+vG59uZVzLfJ/bpXIbbB+I5MuZhov4m82FKml59QQOGu2
oFsbZOP95b1inaPOAE59Wfbxt64K2qVujPUAzqqeFabICvnqEQjTpbzjbBvq11tP
8B1RNlmkhgf/wP6sLmq2Bf/lT9Z5tNY+skdcE42gCSkUit+pghTCyr19tShdkcW6
VMGu2SAVXIhV6D31LG5A8rDR0MmlyAQ3ac8dkfevbwcfVW2wOkJEFamyEIrespEw
8I6IoTLp+6/AYj4CUUZLy7c6UAHaEiV7CGrsvqQGyuMTbJmD7AISmRic0XC94rCv
xyamxEJC0kn7iL3UBeZ4JpieOn5rN6EYQaykhJIpUByteNWurMfu2b9ylxmhUNAp
/Q/25kefwXafP98fJOp0PbqAM7jYe3l9nKLulK8U1N7b7qP0mrPTe2fMxDzOE+nD
cbdFt1UwJFtnhA1kelke0ZIG+R5emETTTneWbtyh8wdjVqgE0veIwuVLyEUOsVQH
anB3Axz1nxbnyqFHsrR8AmRHzLhv44W+Yv0X20ljeRAUfma+WG/eeg893SikNGuN
+kfJt+CSRs1qRhcdX974tRmeH61x2ZVGCWYQPBBIp9+1o2EnVtpOsWLq3roglSh2
mh2H9N4PUdRJDnn3bnn1zzYx7wbonTqLyzuk9H6j+Br7STabYwiDmMEQInZnxQSN
g0JKSNSIY3N0pFqnViwM/vG5lTzljJH0V74hxI+X8D0EQQK+dzZ+rk/OCWGJlZFN
XsZmikcFYTfgqwKFSSR5DN4kIbU7CyP/prsureUhTP7U++CFBbzZ3pSIG8NKu0Bp
dvn26ljDnsLLDPn0bypvDw8TabB0uJFvklAGwGKAF57lBePcROaQtUjgZPAPcIAS
FTR7oeK1gIRQDweTEKUaRUBy8wh7C+MAUXjVCISd5CR+JMOA0w0DMWaxSEtNVO33
gjd/LT2zSl6cRMHxQqZEl74zQ782s6KEyMLRyY8olfMRImfzxZhpcjJBGlWFIbVw
pumLEVmj+H56eFSzZ1Gs1BLZM28SV3sov9ylt+y7cPp0BhYWM+tDhpuwpzLVj8mx
hXl+3aPbkTmCwFMFYAcEDaoRGQbLex5+C4eNzcw4pe+VXUJaMKQQDE3i8UDv3AZO
avdep7kDCgjcoHbPTCV2AvFvneMaUynKFS5m19vysktuZ2Nm+3OMrMQqTQsbcy8J
WqBHOknCKo+KUJ1YTBTymg/m3VUFSzyVVYiyYL/vsPausXB8Oo/lFQyaDa3nBNgI
wC5LkniRx/h1aVB0VVWYjw5Uocp13u7cqs4kwbG4Q2m+KV3z6m3mROyRRUPLX2rg
Cmi3ViQs/arBkn4Rp8ZbvyvCvoqZztyAHdBJ1YuAanZ+VC/GUzPY9KKj+NYaaB6H
fbRfUjXP/TswFksTBKQRVqgUIPfUDOfaYXfX78rw9G/ngO0sk4t3tAZgxw/U9/Mo
sDdVq62uNGNZKJMnyMml+BHeIeDE53XzrenYpbowt8VL4eT/f8GCfFsrIk2edJd9
Tt3hj/hmhWZ8f9ItK1jVgVGe6n8cD56W4+TmqN/ZV7vc5VANIugfYtcdHarvNOgJ
9gH+/OcLWDWSqEanI6pSiuUE3TKQQoMNZvaz/3/ZsUd76HQY5VWWbYiNewjHPmT1
L4AxXSr0XpX4y92fB6xG7JJoCUnKjmg8QLJSxwB0XkWmyDAUhGc8Zrpp8CL5S4mt
AMDz1TWcbbNvutTi7arccqmed3RLZf+rxdA1nxeu3dcySmfXBRox/YIBDJdwx/oF
979hyrfg9z44JtP5yZHKE9pEetUswtvw8SKKeOHpCWKGIY1r+qLK6v2oIVKyb/0/
2oR1KcmC1eRGYEe/AyzXmL3hJGzno9UOrsQ2N9p+ufpHPBi313Y11x6uOZt9RXWH
SuorFRyW184HQkt2xTR0WotrxGpnLRpgPrg5gFDS4vXZJbLjoqzlCYAIOUAYzD9m
G25bPoYJA+/ylch0KuD4Nnmm5eeb9OixzhmVfXQVVLAQl/Kt+Q+5MukgRsDDzSqf
At2LwdM0Mw/U5H0b2AeWrdkGTaTJVSH8FQMheexUEbsRx7iI8q6mVpl0TuCpANMz
sBb6Eej/wqMtAjQx3WAauuDq2h16ABJofl88aW/+/ZsieSx7YfPZJIvYifwr6NCQ
URFPrH6l1g08YrSANIC0/mG4l6aVgI8FpFBxHT7J620O4u8Zk1Fpd5BU0HenOaQ0
3psFc00HNmqAiATBghvtkO6HrPCf1RbU8P3p2L72H7UDLqT4UQPjQDlN6Dzbgal2
GgeceDMMx9eURmVxBwR7YTXcaRqNsUrJGYAuYY5v9vd6dnZ76n0HL0j1LvoyadcG
TsHocvijo0y6XOQqOPaqFxges+lO4AjgVR86/yOgBxzEfzJ9BqbktlQpAJy/qcIo
ygFBwi6QYw2LVZBDWm51pD/xzocpIzPne+cbGI0lwzFXW1msER0gXmw/OsSoX8lc
nhpZ7u3J6CYy43AfJXcObfXbCS+dyNJGt0KO3H6h1fqu0yKRlyCloDj+gsrIR5TF
pA+8ho63aIGjjp3++281LQEPs508jDUOqyPUA0jUex3ajsp3Faa4mo+wMi+t761d
/0gPfuIWU3pnTxhVA8IDyMq0SZNcUurFkGOfJFGNvflhZ3Fvpz5ri5puwUeraiJJ
uUHei0olNwIk7PRxawFOVXXgxZn+tSYQhUayUO4njcoIhlRjQ0dCHAm38bursAJ/
tdSVFsu6w1vWUkv1L1S6cG0i7qIDU7qvXguC7KWXovFGCfzc1O8ZoQUpLO1PRfsK
egM8zmAaDFh3bzcZOpc27rLogaOnheJzVQfHEKBApoaFyro6/YC4pMXZaJbtNAON
s/nryl6QKPfKhsMwCZCFGBfY0kBKFFQfONM0rvxKbBNdMDu6y4uPlY18UvtmOu+/
tW9nbAfuQ2ORH50iEU83zUh8QTvl8YkxQTjcm1DmYL/AR39CNZDz7eR5z5+jvpMt
bkI8J5OFmuAAOexFBnwzK4s760Ym7xXN0r4uevzYn2vdRTs2+aZqSeicBWtBlzOE
/0D6zbXCZ4H1nQdEhOfeRjTgFdg9x2lTNXTWaxGB63bR8peIH+0LgZfW9R5xYL3d
U0yi5eI096WSSwKg4EApzSfND5pilPHfsqDkupl6jIDh5+y3Xz484FPHtFpXlsG1
nDjQLNjP9aB58p8q0yTimqLMHc03F3uSbgUARCthnnxHITfi/N8ot5a7w5lhXAj4
Ww7G648VxPfx41+Qd0lcsIYjLFzEehr12/GH/sr1gNJgGy6OyTqyZiBoFBDqE+oS
0soskXeVdlbDjRJm41X/1W9kj+DHqJ2i4AtT7jbd6cQNkV0V86dZQWuqfjJRhFid
fdMS0vHj64QS6sn67WDlG00VubIz7H0E2AhOQOHGZP5WFsE/70NjinUPQC0z7SIt
Q+PPCDDmnmWsRozvvhuOv6njWFh2azCoM4i+TCdRDCBbV6R1U4vGkKXoFYF+9HKl
nsTVDDXCyWtMeE6E8y6/NcZ9FjhT+H7TR5LxiNvkOguPZsUs6+RQ1f+N7oloXfXj
TvC1PrsWMuJVMnvJapus9kPOdpOSiZLHm8nkBTsvF6l35tWmbi3e7X6TmU++2ngr
d7SwOIvF2O5X0tjwfiUzOgeA+NWWEfP1+g8BRoLhqyEyusBM5Vh9IgksmQuVQGj/
dDUccRjXo48FU927ZmeQSlSKjih1Eo8duNUGKHbLFxfCJzsBHNBIiOrWPZS4L+v6
GyhRCV98wAZDJWaD/a9+wlRvQTwgQZUU+1+hrebMAw9V06cWZZULRqTrHttKsYQr
qYOxrb6c0c8FsU5xSYEwyYY5CtczKb18eYa7zYu70Uzwsf5SvOaHpyBXHIkcNwlt
dCSYE6Z3RXpxINrIPUHBEb+eP2A3C5NhebLcWhVqI/bxSINwEev8VwDZWESeu0sl
AsPvmA4XhcDBuCSw3nTh3Ga9kBKJ1CtGLKoyCFvWp6yV337rvHFdsMsz4zDD54ko
Eua4R9BW4P/P1VHu2uHKqkX+B8Sf/UXjemzVicyUx7XRR+91BixmyNzDJyed14zN
9p/LHmO++05FXOhadjR1eYBPW17qEKG1ifpNniOpoyxGU5JiKJgx4N3+kiM/KI9O
c3oW7qX0pxS6SEaHhXgUS/BjBQ8kIsNHuMSvKrkeBTbjF2vUVxIER0lnZ0YNUBrf
wILnDWk2gtbaUJSDl0iCQEzt8/oQlgFin2yl48dUS+JdmhKMpzBJgb38Hj4+Cml+
1aEWnhT0fK1eZGabTqcnW/lQ++/mmDj9tE9H8yomlp06Np5J3Y8OAxyvcxCVTlJv
nhRhyfAjWPNa8aH9TvFZHwseXPpr3H+FMdpi7hYAZZYsx8tacAKNkdTS5glepp4H
/bwfoDBkoM0zJrXsQhal9w4DdwWXC8asfMnmd2QdIL9sq1FIj+n75qta95gM7XFx
kxXHZPhxLaNTJO9eeelc467GXa+f6SMSvxQ2S9Nsnqyjt0W6udLz+3st5WrIPcvR
sz4Kb6HDJkyDTbWDwEolkynisr6PeWsYtsd6Mkl0ivKuA3JKJr1jwRmpwEX/38nJ
k8jULuGIpEnkO33dDNDtiCJR8S9mxnBKHXlo+gouc9NjhxacN6icoxuFqmubjbJy
sRUEo97r9d8hjx6kSA9FzTWN3GtAOOIeA4FvbApdrj82FCrWCBDbNJ24UnrAQ0J5
vBvU096OgOyPqHlJLHM+x4huRsOR6dPTje85TxJ0Kvq+2mKRp6LVJMr1K/InJEam
E1VuleBnCqt7nuz/pr7JUCa6yPMYIZxhDRu1H4H9LG0bms8U99aw9KqB02/Clqj6
bMFFpALUm+I3PFLQRx15eOmFzxSAH93PEj22F545WcTmvHtu1h6YBgaDne3HENcS
n1Ho4pnavWD2+15fRNzDV81nNMFn6gvolpg9TEAJ/aWYRVsdgta9sAbDOHoAx6kM
lcEl2UfQ+RG71QUK4su4cYiYr0nYzNyAgYFhi11kWbomtdPnXAbZnfl3i4zijAKp
5Z29HBsuuJQXer4qDMrxlJxIsCY3tTjt2IbvQiPGckoIh5J3IZwXq946IWi4eo+r
rFgVl26HrIFdO2jItCY3IryBHahJCG8Ep7kZUyXXdOKwvBP768PIVMVci4UfhN6p
9L4jyKmLhIM6iJxlrhPrB3nx6JU31YXnIJoHvXy50yXCjZa7srli/bF6eLnmY2M1
2BVwunVK/+S8p529s/2NwRW6MLzuydnTizvrw8l/fs+iZzkCzFuFIJ35Ehj/g8Nn
2eoxbCkNmUY2AiFp/oLwWTO0wLARj4gkMYoDWC/X3WQHvZTTPMaZX82XiFZuXcz3
Wbkfvs7WBPp3Wj932T9IvTu5oXe3WhwiVpEJKdcX6fSALKSqp+HNYrB9q/GDSX/T
yIxQ4d2I2bt0f6jMrsXQqmvs6wmj4ESbGPuOLpwvIVA6Akd2qE4NgPIOXHUovN7C
FZfCi+WpLJRMnROeYVPbBS28UID2dT9+yaAbL1TOJr0xkAay81QKjevYK7v2eUKm
n6aqS+KPh0LmwSIPcQ35JKAbcl/guk8Qoe3CVamqGFHxKYeItd3il7bUtodNOKNe
RzAjuz5YRrsyz/ZPpIhjpbB5P8mvJ6HlU3OE5IqOrhZgE5C97khhMPCKkImAcpDI
iH2JzTaUaja6ImjWZL4LO5SZ2b0eW3/xuMsL9BKGtdBWqdN2TtYbFd+CI4kPn+UP
wP4rUBR94vZHW5uLXJBzCptgXlAdkJGL67bNIhPNeU2c6WfEivAsshHctQTO32P0
AzmASXVozRM5RwmDNfTUvhmYZjPMLQUxiBMpcHIiLjRD3n/I8a4Pqy+wcrOIFnBP
a6GY8oiOm5nZSm16gYygJ8xLqjei5hVAQ1PFEC7ZitFBYahFRnGCPfg5qfzRSxad
Co+Cij/wXfBvGAFrWaYTD8G1Mzslq+JG1swSCCuBqCVB5xngA05qRdhBgR1BBzra
VN+zHJ0gPe5++YQCQcDop+K0l+PI40OTfofpmEP5v81fC6UuzKtaxt3ZVmACkXx3
VFEW454jOW+oXfBnr97lK0yLOjQ44AtohaLnyj0XtCT8tHagHtVPD3lXY7dKP0BW
m+KKOEpERvT5cOchmVAcKYpIcziW5X+mPOYV4GdgaAriayqcMJvIjg/SHLTvX3g6
kr0zZOT301qojFQijB7kbnkBOJCglFBYSCSKigWm0x64E0rIUkg17xnW7qsWRit8
kkVUHlfWj89dFI0wDoQfpjuJla4y0SlPXOh/BESWPBF0zS6Kmm/aQu/R5oS478w+
tZ3lLWmm2ujUfm+BbZ7gjEUkIeGvCNM08RiZyHdc9ZtpW97NBOMKkOvzNsew6caA
yuB6H634kOcVPegHg7sop9pXXxBnWJ3oD6vhCrWi+Dt0yZC4F1GMJVavq694fCNz
djIsBILonyJq4jFr16+P68YIIG1WuXcW/IGbuJHkjm/8/hvr/eYlDMsYRVbUa4d2
YETjH7m70IEc0kbV/+nodZAxuZaXhGnBEfb9QRxfvOEEtD6yHE00cjmVSmR0x2ys
SjYSs2VEpEDQlQh98UtvPnucAi5FWTEg2+VKjYYBYAe2NhauNrXpEXBUcqe7FmcZ
pQHt/kw3HGWGrRdIWoJ9aOObZzJ87TwfMh/tXN/gwShhpWppmDnhXD3EQW7SKOh5
WivGJBiIL7ZjDnD0Znptf0W0yaYHtKQfyVjJsk8w2fjKV0h4rTQ+pSFrIR+jgSgz
L2PPU9RpYxrQ604Oy8lybTt1qyij2CHX10zFeneo12Vp0Ap0SP1CbP7kF96mVKez
tdmtrJjGFxlroETLUX/Yt6g65nGWNUu0VZGKh5lYWVh0PMFqmGOqJyWDY3eEC7Pa
/sor/mQR7PR3XFEwW9H6KgvuPFMa96y9aoGHfhy7whfhct+tvHxHvHvui9IiJx/6
zsso5vuXk6xa+g5O/0T7kAdIB+FClVjTAU+szX0vrIwBtInpePWXrkhoEAth2DHW
kNrLxKG0ylVg85qj6rBjV9MFZoqdmj8D9jxS2deOplMmgvwo8BlTonNGrUPWvTOC
qUYVZZuG6mUkDZwYMXLmIGIYUoeC4Ufc1kC/7tdpe7sssl0Nps/bfWMvYfs6jBPi
ixUKyny9df5HvXNDHcAi/uGhg1WDQpflW1eWJQBmpKpHoLPnluSs6a9x2+qnt5DB
FKkFG7o7gKuhhi9JNaJWOg==
`protect end_protected