`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 21376 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eislOGByxcl/gRn8UziAa+H
mjgbsd36EQO5Ail/O6Xu+Xx/ROMSlvuBazdeHDaf8f7LCs9GQxL8P6focTE80jrl
6rOPdHuvc8qPoi2M563aKcF+GDWDr22cj3ooWEx7WV56ernDQ+XwgMT3+rJT13jO
3OKzLFuXcBcA/XRAU8EiBVtzwVoqxWUYvyJu3KbOEDBw8+iXyqCT4yWNs2NgoiC5
blWJ73jpaq+9yzw4AWmT0GF+SCqON+xjZv++zzefonb+NXVS/uuxCHFx6AcQII1X
qsjNHAqNcjHcTt0VNNnxQz3+FXnJZLDqzrwnr/4lI6qfJiolJ4anBxGphlm1WKWr
oIERMW3BYKdCU8DtOHWZBaD8cDw8sA6/p/Nc8bOrBjugvqCQwpIE3TM/ikt6J++l
FzbyOAv7nYR9VupqBpM+jBXdFF6GVOd/aDPEJVz+Bsi4zfPLmPxgDAfX2o9WO87z
pWENU7dMlMFY2OUMiDxdsjyDUV0+T6/MAKI8Yh86FVsAYNcRoxMg/M++1NfiSUJq
15+IyobmWTDoEIEQGDUKnuAnJi38m0DmqSmSNYx33n32Luffra+tX4vZLC47/sE7
OwK3QqhAvt5Pq9l1iknQsRbdIrza59HMUc0crtndwQrLQN/pQvWHazqc20rGo/Yu
O26ccbCoauZa3yvpz9GCDV6jhWBKujKouFT78wQYpyN+8M5YbirJ83Tdewid9DfB
g02ppZrtp3v1qg4QAb+F7ByBFUOS3sGtz8UQmIMcTEavDE4Ye7FWf9VBtGePwNhu
WzBm8jhYqSoM2kDh1B5M8D41lcmq0AtdBxt0yajPJvfPNGfKBSF24IDwXQFdFTE4
D5iUkD2ky76mekzi7aIRC4h91pZlsL2RRRJh0S5PCjdAR8f2tBT1lqOg1Hilbm0Z
WWmbvq+bi+tRLOxnfVD34D/It/7S9fCCC4CHJZQl9Y9Aow7SZ+5Ff0xrEjTKmgWB
aRJKvu5gmm7W3VWx5yqrOBRlB7RFk1EP1tT9tCCeHax2kMkBQ25RclRZoWHZkdfY
ZKcAHH3h+QGmSmhLDt80aCKe4Lwre7qVNIlh9gyfkslfh+smMLY2ChhF0OXUAdwr
WrF8zmZ0ObBgYFV1tUAJUvhgQBHzcMw9yplMyeHmbHteWGMSuVxuOgyPrg/AeQ/+
nf9BHfu4lS4uwPuZQBi47XPKq/pRGSA7sva+ZOXj2nnF86KoH3sXj/43DOWaCNHs
E4mY3SD6RLpokFqJTaNkX+sn4FdFJpsceqqtZxWjBPeiD0EZ10FNBmbMl42xD8Zn
DzSTqkqh5Cnva7Bayg4CNLVxNOuDz6faEQg+mwHtKrm4coT+e8bi8djLy7dK3Gyc
drpBqzIfrQHmK0vuSD/FwjfL4iIKA7Ec+e4/ziVm6umLRIrt1sJU5MxcAUmd35vg
OaAa6Nt+xXEde62EOJrY0sJBvnSS4C0guLs798YtL9mA6UEf5Fssl/qXkTiTRUX0
kfT3lI9sgDXzBpKVwe1v3lzPS622JOk4eAiG1I7TEp3sZgcgTWQPBWH+A7eHIBEp
1NiBoL2l0pjvxUKroh4s32phS1k0HrKCpXN4hbizPtPyh4TQNIoC34yRD0tw4/6t
S668gZmU4o4LELDGzt4X5ED39ch08jIfUV4OET+9bmGEippT9qTayhnCxugJJ/fm
xx9hTlDrt686F8lmB5wPGSPiXz3IeQqOY1z3W43GHDDSE2JFK+Gpt0P7CMuCvYuV
3o1sUcQcuKaKOdAJxc+76xfUKiqVjsLAiangbDnifusd2aN1ytDFMpUdaknUVlP7
vUHplwxuiAD6IfOfZMYmecRZtW4v29PRSfTK5mHxoGBi4qiSd7OzxwvAX6nNyr5U
rXorLPOiE1Eu2SOpfv9BfYt07NYoy9hH6ESO6AZyf34sePQACpn/I3eDhFtGT6vr
VhW5nqZM4PYvOivoc4+pU05om9ipQrc5V4FUtNUr066d4Y2pfHsTpzW0G7Wn234A
a2TnRLtuRdtfCCHHr8UXPmfgxC+7tkHC0/r1AxKt9VRW+oviU6Zt3n8YL00W1O4l
7D6BGtasnJxwWdnyf/i48WvPUJLy1UXNto9GSEupTTs4yGNbWYW8Qg+fKVjxboWO
23sSk9c1TemcjyMyMX92L9uWhSvdH85Rw/dPtNKsH+rdUf6M/70Yfjhy7qOgNxCT
+j/DKP5f6wDQg7fbpfNe2CkkjTdU5swag2V35PVWS7eMIxZV1kiScH2bvBvwd0aS
hWQHfHubSYF19JQIjv3A8kZPRbxpBFmu20NghjWyOW2TtFM6mEVzQN1xyr34hvzk
RGZJOBznOWlIZY9PfP294YROAg6HyTOLHhf+DE3m+zgqv9cRzXDTVoWt/BDsx/Ku
DzUkL2yBLqOgKBIrz194tkv4/lf8Niu54QqLcs8GGCfHGWLtF3fvRuEjRoSRgYPV
MOvI/JBBhKZ5ugGUrlqcLTmdq6DSBERLaYrdz2vbyUgJxR9sZ1ZKlIi9MCz9QZwp
+ubEQcQVIE08366zoCjhAKovoLuOV2c4BI3Wru3lfUIeymvpL3iRRs1l0lrK/IGN
pHvtg0cDKdP1ih4EUj6Y0gqKcj++NQxiDoZwRx9SRpqdFwCVyxfs7FBdIUg6It44
kkQZPadUcbBCqfbOBMlq0pV50kiEywS6MTwf3I1PAofucbgQ3PKR7lbUS8n2b6xK
hFc1xXvgscdqTnJoaVNQA3doaMtN0z0dqPBDm8aIh2rGJ0gWhEPOxk4eNNOciESq
f9ppwjYILhFEMA8UlxkUytycatCWXBCaBTY86qvgSysCOvPUR/ycg3EzsZHUxpVx
gINNFGniB3QlwOBdh9IEbMPp1RKKGmS3KzJVOIR4on6mA9pyk4ULewpbG+qacig2
SMkZGgswhHenOPle6+4jifVWAHzEEtbY1KHCVGbcoJBNWMROIMsrQVMdF3/Y7PgV
hUQoFrFF8VtU//L7Apw9/lY+YkkHXqN5EOrFE6WonKtnth5Lsn3K0WP2SknZwlTp
9NGi2yZYf0Mifszmiu982QvCjonrXXg4QezfCJpceVRedhME9DYe3yPFp3Q0vMJ7
ukd69QqID8S1Vj3o9DwWODgTm8ILjnc3sDwdYH4LkxQJ53PfMgq7zuB9Cf0p6SAo
ySy4j9U5xHQM/7LZFqlWn/cCX/Wby0Pw59VdToV+nMCjb3pUxGO1f2LuA9wUu5Va
jhppy/0pIoJ1VDUoOI+JlWnPaUUsjuwmFF2Jjfy/lem37d0lUJbU6KGfEIt1jWoS
GLTERIIyD5GGT57DQKGaxLzjGXHJR1twNJRi5aBG8PCwKrLPwicrMh8TNXmOsWom
Cv0NkioBU5w7Sr67MBeBnqswPX71ggtOhQUGBGOqxkNkC7z5j8Rl4ebr+qCQzl0D
TKkveP1YyIqVSxit7WRDQo345LFIyLXXKGvAQ+A8rSk5w8pAXR1clPfIxhtNZ6nU
KZ49PPZl1XzDc1+Q+czA6RMTxmXTbe1OZ5GwXIV4Dd288G7HfMgOmmIX1dEOssuv
pMCcHztMy8ujiX+4Ch8ksx7Dh4xUFvW19/2H8JIxh9QVF8z9jGIvtcXyisZplgg7
ETAhpJ5PSavL8ibWeQL8CAWZDdJkp7r8e4WkUYVpwebSWNZpSmbF/hj8r7OGbi/C
rNJwHtiyr2pqRf7saJmm47trLyhsXeoWD2xyIgN0lmgizRc9awckHg9wTxDCcLE6
3oxMT3tP/Xz4uDd45f4uglaqjFFm9VbHEWfw1qjzmEJasVLUQxn4SBDUIfvYIbqu
RU7dXnSz5cSphwIMR3qfR5e70yc5h0JPrHSn84n9rYqkV56HV+qHNvqCo0OdMlVJ
Bph78cYoSPvLF9Y+ZuxYxqaj4PL3NFw2FlIiA17DWlLMx4JmDvZOVLMsEXLfCO9c
DXwEmUN/iKST+WBptelXid8Op+5T9qK011IQwsKIioBiNjtAvwGKxCLhJNF/IBBl
KgopVuI1SwOW2rAWWSclsbvqlWndhw1lM60TkWauQnsKpwLOYUP2xx/BRuH9utWB
u4LcvsE2ynaUOxhVRu0bRBt704DNSJJ6X1Xt4ATDYT386fqGXQ0GKXAJ2m7yDguT
tqg09ANkvenHJqDHVl2+4/eXvxUWDaRAHVMPMrgzfdIutw5CFra8Mg0TmuglfcIR
38JJNysda56WeW3/D0Zam4msks9T4fOADvX+LE+5/fZX/jf4ukAmEI/5422fi/eX
7R9XlXU1PVz9YBtSrp5nVVDT9QzXdtgwE7jY0x9YyAXt/XZQHBuMjgSugVBpWaqz
NgUAp/p658q6B8XS9spmE1Gj8WQpHkQTBshdGQfEnIK+DQwqLhJMHX85tyfXn7Ap
R1eluBUXuPvindajBIVhfaENm8aJcysR7GsP7Se4ign9Vs930wt2HGp5Ec1BYXPL
htWhZjXJolJ9xv1NJ88hBbNoIpxkqWjy/sIxT/IJnxQ5e6ONDs3et5q36beg0gei
P4IkEhH1kl8W8eaOoGdTz3G5VdkBM4Y0zPf4XOFGzrODBECJnCSX4XM6GFmTbrS7
B20lH6grVey3VA8tq3G+yVdPBZDUiBFrR+/ae0HGl3YOHEvfIVLMfJDFrPEUmNh+
aShvaYtr/ZkRYe8CvDz+5qbN6wHfXvwtj9pYQoj+luLfqiP+GxRl50AHjHdbvMD+
rR0ikx1j8QSVXTGrKwBGDZzLcRE4JoaIldeabsHcNCjwyYUqFR8S6im4ZrdY2G1Q
6ij51unzYe8qaITOWhQUnqHvVJIpmN7l4pcfSqyCe+omI5mA2/O+HEZjK/V5nqxF
ovSdTvMa6BfWY28DqFbJlOK7fDeTbF6Na8pIBezqJDUc6hvFn+k6miYAnb+RXkrR
+l8IsSV2vkn+qX2ySCYgI7dTc3Qp81l0Jo+GlDjHTmVaT0tCHUwklzBRaAlJPfSM
KkyXUmCP7gpL2AQJhA72mQ86DS0AMjGu/5ySMe9wao74jsYyc4sTYHCO6CLmhVVk
5IHwI5gZ6VGKYyYfLn7x94MtbBqj6SvzJ1oxblA/xLppEKXntv9kaCpMkvFvTHRZ
5wGOumDV4cCD8SBmHkoDK3acNbFbf6wyTcbx21ixMA90bO0SknVl7X/P7Bpb+t1P
hLyLjzmyxRk5vzuoQQe3c9eEEfwlR+zio+kdN2i8erT8fHcKE62MipvyXmOMHexN
t2AWPipZqzNDfX7fGf44RAhfTiFg1BsE1hQGBMlS6UnLQWcacr4lSR1qhZNxMvSK
UF73kv9L787lhuKFvYsKU6aIV/zWKQJgZZ9CLo4aYmdS34T4JOmCi8Vc14kzaEad
dYBe19UOgm7C6BHJnpL2JqQxQCQ2pB8OIl+ItzPaWINLBVJiYHjMIWLy5Q4HrjGt
FBnuxvP7ZtlppiwQt73cF2PmXbLut6YKTH07A/fYE9kt/bVSVLk5F45Z/EKUrc+O
TE501DQawSTE+DmgR71OWA0zQtX7/Fov7nrntefVQ8By/GDWaNBhDCKzIrRQIs1V
9jcSJDa9m5qTco3/z0VEOD2edIBpKXN7Uvkp1ChKk7Wl9Tl+qgWFkHtN9tTEJr7j
Xr0B/bz/kcg4C0MwpJa2tkK98tx/YsRTIlAIMItlZ4onj8pABkVrvPNeRGSfKc7t
/2DaalIOjGR9+onrUNsCyVVr/KowsN4UW6AJpI+1u2XfYoEOEUG58On3T8y6GwYJ
hJ3dpXqDhOGA+vOQTroEO8D6mzwzR39ZuPWmPcJ6HmcEzBIHWX9Ymi+xI5I/ALOs
W5Hgx4o4itNoQWUuXQQYZtedF6usHHJHnYcMwbC9F4Bc8lDZV3XWVFEUE6OcA14U
yVynxUiva+4DHRtu8qN6XCXQI9e8U546+AX52WPMMVWwxWr5IY7pWkY9KmPQI13Z
/DPjrSxeo0PRSFvAQzOKp4G+E9hApwKR2BBccOv9z7L6pw368ZxIaupBZbGjXzlB
C5s6gFQxEwQ9qPbSyiONQ+L1Uz+LV6+VymwubAoJByX7+COG2xIf7AsSnYlGLpK8
7kehhgjSlP8R3vRBDybYL6TF9TBUL6ameiuYb+wQ2o9tQmMqeY7quzmv/vQUw6k8
ZE+X8dQVArCu2HysNgDq0iG/itQY9X2ExHMKRUY8Ypd/3/lFPlKs9SSuMxpwqD82
hCotHHlVvsBBsujDC9oaygroAra6mzrGkIwW19r+SdXPOxyu3EQ62JMLvYWBCpdf
MvY/hcM1+SlRQD/fkM5v4oLz14UFouinSBZ+7wRiH3cUlEYEQF/msTTsUqcnmcVL
nns76Du5bwD6xmoCSM6R6dV5XBpZvdfi2UceU+hCeZMSNGKVQ5AEUXR7q0l9x83Q
X9x/VFYQtc+GIV3E3rqaaVdGXfo4783fD1rNJuEvANexEeic/S+sIoLHeeMwm6ve
+1HRhbK8WpTSGn5KE1mfE23XDpMXA+Yu23lWfejSaykNdQl4VgQ6wAQDoSXUtJt/
QFdjZJ+irI81Z6DAxpO6c1BL5Tf+n/Zq44lOMeBafKOY1GXe8mW90gbEbnwk7KFB
WDmAWxH4WvO2UTbO50cgrPpUgdkUjEJkSR30Yktc0B8RawDoUjTyq6KZ6UeViv9T
ekQ4AzITewjmFjgm+5Qj1TGnyySHwvLGxEZB2LJ4pTMDhJ/ovC3TiGJ07RCzAGUV
h8jxNE2mzfI0K+ADTSJgmLqDGCLBqFws8LRXIPGzxniZXDO3uvy3Bg4zyoHtDrdU
8bSXz8iUv2vbbu4eJ6h94O0wtyiUTbExeHv+I1CvvJtVGsr+7V7E20d2bQL3RY8g
YRKwkFftdGap+AW+IiSjQpEyu84CWna7S6ZTRLRRjdi6IkJfcHzsGkVJ/dPxpaqT
bfYX/qFgbmZLEsM45slUGm0WPr5yu2RV3bQboXvt4aCz/CWzptlIOhPbXbHw+E8f
oQDhoAxVK0ro2N4W1wjfGZwhlNoiQZ4wTjvSxC92Che1xKURjqxQZ0ZnJ6J2jS4Y
1Ro2HrENc2eaAoHwgd0kx2D+UCIKrFEy2Ec02vDNumxqjIGqy86VkvVgI7mShKq5
fj6wxfHiFo4KyD2m4K8eow3+JRDbtU1gZ4uosfy/eEZkgBuvcCOY0vzIBul+Fb1Q
SzxMLtLFMPfp1ZIeB2XhCy+KXeisbkDCPQ2ZtHGxENbkkycJkgpycotRW2LnAc4L
VUDqgJ3dCToVx9rW9GPbYtOnUFSeNjlejHMlGK1Drlv1pwAgqnQ2wpnGWFYsePyD
KmWoyc6SrK4KHUe3/0G5C9GBMRNOSRiH8JQxTsa9foc6t8zjXm6pQJZBC/6gzuPi
0mx49mYSt1G9Wk0tyFzi0y76eAaBJJ+KrwDAXAIpzjY9LzwDhQO7ohgHfqXyUIi2
AI3WVnOXf1vCm7K7QIG28JRXUbu6UUISFZ+2zodQBmJ+UWJu42lrGU3b47chauiq
iuShzi08LhCA0qsovj3b3+g0XL1ja2u7xPuKX8y+Ghwv+moIw2InggEzzyn0balV
8DK9D/jSRQf4tHpBHAYcqqxlB2iNh5s2Dhm2SZ815Acf66Ol70RFngMYJiNz860N
EkSoFCZvDQM9YQsm5xAecCAmzgjUIkgnBGCXR208xCp+unOqlU8ywW9O3JZFhrxb
gY/8wvv39nctwcEBQQ3xYnq0SXxXYvBl72wISmwg0egDmiQYp+WLUrTZlSMsxkGh
vsdQ9Xl/5L5v6kEy0DZZXKnvENZhZbfIvzxYkSfLJiILjVzOUFNA+zOg5o1ja8iS
HZUQ6Xcsw/kQmExwQyZi/7zfpSWtlR+djDIim3aYt4W96pD/sptHkC7P9fxtBFm+
k3CZn4lImRsPV3muC5KEBzEOaugncMPlCC0AhXktfW8B6doCsYZf1KodBLGWYUj9
xY9Nd41PHYwQp6bqGmjfMUX62tCA5QqSy7QpGucs96M0ZhP9WUmpLdOTplGTLxic
W4il+ZdzZVxtv0jLS5CeCXfmFgAqHpLKnoqINQKtN/vzU5PXyVHWq2rcVaj9iivX
HPP1uI4m8YF6iWilbOyZW4GtRNSHFdM6KSbLgQcqWa15b5j7eP7Voi3oUna6a7rT
Lh+opbGvS709SlyZNBGkfkkfhIa7p7119sNcf1e9nSDJ2Dd+CIn4RuMFkogxZ7nt
uBZZWGXUoR70VE9qLrIl1DGfdBvJ/jxjGSODCdXmkagBaCXD3eurQ9grgkG13/57
jLYYHS9SKCmlutDD9elVsg26DCMlQAFCDn8cXsI0oqWtof61jeDbLkGt3a3ZYuHz
u8AMtur/lx24PpdiEljRTU3xi1AKfh5o/Px8UphkGFug5UehX/OzbWZmi3NZRlkR
1W/hQCVTBSdBI/lYVxRKPWZu7/MNo/99YMY0DRaFNyf6RjVPRtn4QgH2yruOJTJu
dTVrgYybHyhgSX1+/F1Ac9Qp+d8mZU2yGlkY0kDIFLietxBlSc5+3lz3dLlWq5Wb
fUZFA9cFyN9/JQ2poP4g1NyUwqOLLxDPA+KJn2IO+HLrDVm3iOZE+nJzXqmImnLz
Iri6N70UdExdP1luJFGWYrBxXriJ0p0VsS39QnjVHLOAQwTD5u6rZofTFqSYqIdG
sT9jxrwVei2lBBGERp/CqlDoirsrl+hAL6TQznB1Wtp1WP/TVUao2wowZluNJU48
ZoKEQhb8t7VAus4scCGdwBQqZIeNeaWcsN/b2jZerFmbrt3yMWVmHYKUlZVUIRc+
G45JxwbJuIJ7IAThFTjJ3M4lV/phQ26SZuekUbZ1gVznEzie4WSAZopyfPNwiVje
NV1KdzvLH5aMRXbYS36KxBBcuc2q4dyadW2bVwssc28k7Dxi9mmLR8TCtBLmceN6
lftC2yeigIWRPRfrPAe042R6U2icOLtaahv2MliITyDxc3vg7zJT3IiR0lvau+Q6
F+2+rurWl+A6agbxZf8niKiRZKXHkjATnAKPQEEN6TJWv6FtWLyly1YMjnC460Ff
ukuTiLU9M4u97ZOUbyZCJvXGz0JWG+6q234drTOxrhOyvdsN22VJwzvwgZ01QoMl
pjYdtqP75ZC6DA+Jpr2Zu0RVUXVD2m/okbt9XAGCow8nwT3JGs0BBfCW8LpV0nY6
7IpsDt2s2t96Dgr2ZhHRKJV48mI1WsoMw8rm8mlufnMsuxynCSshJxaFsd2fcL5l
iAx21knW+YsDZLU4qkabI4NHu+lB084yIpXJF96vIUK2TinZJqcYLq7wD2FfYIfR
TnDkMIDBnpO201/E9Fo+7ABB6tODtAllXvscr1azTPlLIW6v2pa7EnwQaP/3doGe
l2MYIcPe0aIverYvkRZi46ZnUcjr6UaD6F1dO/9d6rB0hyyQ35RK6HERiboRmns4
mMEABfa6Dq/C/unuXXBIP0er1OLTHcWgDtvLu3a2qYIM/9LuonyCnxqREtLITl4t
ruD7QiaJEKNuFfXDiaMuiHcP/MhDyewYrx0sAqaRHINoC2u8ejvDOB0QP/n9T8/7
I40odqVkuGLwygZgUdc3ACSP3QXOkeyF1OtezePi7HzS0bY8/EpMK85c/L9WK6OH
cP7vC1gstB7xI0PeaPCnyCq5Bxg9ii/f46kCO0lmuKRPKdPTtA2mQZ64ZSsmilaS
ARBIinZIMl0LYb2g7V032Sx2wgLU/eYC8WviiLe20TFHvsr8wXWm7gpoEhRD0Ol0
IYZxN0VTqCxT4x6PLo6Fe0i7ts/waZzJc11C/QVHUn8BURuSQeq+G4V6HM/sdLZk
8P7c/+svgG/hPwqzdQMAL0P1rdt4lu5i3Vsf+nyH7OT2xxH4opkEYiSKWUoZXj4g
gw5kQxeek/JNPN8wjjVdpFJmxb+66GWIWUf1pycXL9xvG5pAdCIwMsA22mMobWLF
OW0k4oWTyNZXBXUzNcfhnn4ek9eEgiQwT9rdY2mNdNW+BQ2cUKdHAzpLJZbRS60Y
iny9ow2pEripd/JUcoR3niUow5cByR5PyKIGgEyLeUUskP9/n4226QeE+s/X5oo6
49Lvgozr4PIO1HcMZFObyaNGPgT3+eQKMNyAYibNE2ERfHYalNb+i0Ngyy3Z9vzO
6NdyQPKcZ0Nu4YDvGf0lqgWVq1QrgJXQ9iad+nV8GIMZu/ZP+4Y95y4wgM0D/Mb1
wwItAp9bG9oIfcKBS7MUxQ5Ho7loVLJf/RMMPqKZpBxtlwdkIYXV0AO4j1SXE5Hg
lyK+F6aXQxvvQUWOd13TT+StMxleZ8tFbQcpJeoCh12sTKDaeHEZNKsD7thu56qm
K/HRxC28YVJRRv8+oe9IitXUbyNiegeEdHFljr+qlHsOhqMfK9OAXIy6RzuF2AbB
pji5qmrjTjCLnZZ0ddGp4bqQyXL/wqxlE0GPle0sOUWTzxF8g5llQPPDApNsETB9
rpxjqaE3ZzvjhjA6feLUfmmAvwEqL6OeSLoV2Q78siaxHcNWReAnuop3TtrzHHoU
6Iz58BcU0vFL2rKtTQC2gQoc4fKImS/iq54R7BTjea6up+5bST1E2MAyLJI/YYFZ
b7pkICpo54v7yj9VGA/DxCWqHPCDgaPqS3YvgtJCZecAfhkCMQqWltE1AROc607i
5hisDrfw/AJ50Lrx7J1UBAJlT/If+K1HWDBGCqFbRKUn95KrlIRA1H9n5ebyMEcR
th/ueSgVkK3OV0AI5dGTc7ouwBKeg5lVYu+8boR2Dum3oLYszvu6gsiIstWyuTbp
E9Gb9wvgQNP2dOUKKUy71j1986vYliSRsrUfqiZomPr0UYCjcS5FNXR60ZY84ujb
45Nu+yHEHTOMhHHCCqEwRqNX+m1/Y5ikuBNMNuWVHGqepQKb7qKZnNlSqjYvnB2M
7FVO9g60qK2bLMLu+t2Saj9Zlvp+1gix62A/81Dw4+4GVCyd1HDAeaL6MRVGqlel
PoDc/dbixERznfN6zPT9zqETZ2DxsphS/jkusGF8/o7LLG2SSIUdSIADkeH5NOSg
jlsQwWj84TWfJC147ZJTOVPNKHcK62puhP74Xlew0rOiQq6U71+Qas5xVXpSMa84
htfIa81+5KMfbxDHJ0QhQn1HNIsf1tD0GUbpdJg+NuueHO2k7zVmAEfE+ALZW8XB
gkktd/UveLpgNAemII4lTjZK8cyixYShEE6wH/GbX6oYa4RalBRinwNQp4OS+Wst
S7lH1lZwhLQyId5CGoNwKPh6c7LV8o6bmWWmaj91H5hKP+y3czAdpdS/tJp1roCB
G1C0yPQu9wetfFq1Xm7jBKeOSI6RfWyMP2qIZW6UBIPlmTSmZlOlPAZDoIJ2VcYO
2YiF8zkzosEHLZKb93RtVpJ2HYhvqgAW+P8xpYTUKYeJkedrCaBYwrkdDD8kIjd2
vZou5ZT2ojAG0Wpcr47w+Wk1PLCTyq9pibdHKCJm3uQVgMGBwRGNx46FJQ8HGA7K
vdIbSmPAOlrYGtx+MZhnjRWcNo7MGYPj3ENuX0G8qize5D4xQTEe9WQHlPbshxCr
vczDBFSfbVZLNVKJd2YlAfj0s4lEB+em+ELa6+z3bF6hbmZEC6XRCn9FU759UYUj
f7IahhTNXu7OtEItplWx9OdO+xOvz6tHvOKp7fUwb04ijTGNmS2CPl3njdO0oMku
0rIBAEvzy4t8xGlMlZSAyLiU8Ptlj3hWPlHT3roKdt5T/AP110ce3EV7ZMKv9NPr
w5nMqGHWt3lG6CXBN+i3OguYf08dRn9eIROgVki5diTNqBg/olamcrLibfmeteJf
r9EXKzSuaH9qLlZrgvz0+tfxNw5LtP3IkylBtiYMv2RAN+8tZh0KBAaGgWlbkrm5
ZgrRVzKsWIh+TVZ1cXg9nw+wtY/QFvI7xsuoPr1fPmMfJQqS8MDWBJlWQrRNVFyE
qel6jCKQB9t4OPp+belyGa4n3kVnAR4amq89KOZzi1z2d5ka+IVpV0ZtOsVf4uge
NDklNnhByXgsNEAL7u9bBFCpyDY8+R9R3N4jNKJ3PWhyp1v52PsYzTm2jnfJGLuF
HdLLH0Ln7zOHtk7eudrLtQTsZiavC7hlenxRuiZ7kauSCCIE4H9ntzaixrMgBhP3
A/jWRh18t351N0LKImzTCHww0PuSmZc8+0QW0dSAJFAhXnX3QF2b1/JKL8JOx8vW
xq6X2h+8xIvqmyUOy2zsuKyJ4I/9HKzicJLJaPuEfbXVmEt+r+hMP4IVe2DPtaXW
gJxZ3j6CGIBBv8R6sEURC0wpBOpAwuXQlygkEee/DZexy6G8EBzC44dUMYc9OFWx
x8qN1z3SN62T+Q0SrOqTGSrdfEAUkUCaEUAxW3D7qN1VgGFmBvUyaXVC7dCA9cJT
vUnmkRXGZWdO1sCwk/rXYGi3TzmqHSP39xhXyVVADQqDx1yY9CnfWO/duTisqlHt
Ciw20ICkFbGAwNKlPFp8t7ZDBIFy65xKIBvXeWvVYOety9Clu0nVMPYXr501TIc8
1Ld3dqE7HBGCXHtozpfjbzAbgrDZrq0TMD2huvGBFQ9IlekYNFotJ9FQs83t9MAZ
akGe7ScrbyfmyqtNZM4lepH9CH3DZ2C5i2Uoz/BYYXYGJypjKnFpjUXTv2fmCalm
3Rrb+0eoJ0CCQzOL1kk29V4NC98C+A4bg+z5EpJpfHfRG8GkPjF28pnOwvCZd7Qx
aKumwsZJ9lHzPGIyEa5GS5/bTKLRMl5/XKE7AawfkAWXxgjjy4XSadukIspsYuew
7BY47Iq+qliyj8xsqEv0UqGvMOPAkQjyv7RkYdaJ1b828FO4vDeCRnyxY9+DE3hB
QRXkh2QPlL+hOms3F/ro8j8DVvIOqvnQGbpd6b8YdhfCjEz3m4gNIQIV6aKofXVY
wUutCd8hC/e1tvyiu4AO9iZhlladvjNQ2bPfMNffyXM1kzucoOe3nhHhQ0veWOuY
gP1ixH+6MAlAl1k9LMBeEFzsnQ+JNAD97Ds5gqyfMoKVeGwsfsSChmqZDBuLi+Mh
vwdSUoNXSpUFzBA1ejLvG+Zu+3GyTzOcqCTK8W4B6QHyaWG2xbOTktrn4SFXokBy
tKBuHfT4urz6CRCnmZVMKo7S12JchOfHnJIIG8ly4hGt0i/vt3mhZ4jW9GkDu2WM
dAVj5MxrRRY3U9IVVk+gauMMaY5Zi1OKfnMoVPTVzeYFJjwi2HbVZcOoipAJka1t
14riNCqE4QFGASjut+0AXB7+lyC8qeiauMq/rK28ovzvRIjxD0BdZxtadgPnRdSr
K5AlNWvg+cTETFqH+xHRE/DQIXd+5agMkFECMqCtHkOz+XpU+FaEnuhwqF5CwZFN
Vi/wBI2/bN3DobeFXAFbE127q+1dPX1mLC1upzYqdZHcsUSAAvN0X5hp/zPbZ8/T
Ns/3lPotO9hsq+5+OMmIoNiyRe1BGDv/40FXZsNdPewaLXcHGajvK4cZjVIOyLcM
u5rW+tARpylQ9LzM7HSVTiLveSsrvJJQdsHVZZbPUzay6A/TkFSk7UmuZXC/pu8P
XijCqcO3akUpqh4GnVCet5N1fsukq/kUBY74ppoHHngvfhLCkc+WkryzINMz49Sg
/xzGT1+Pf5xbyXv1KmZ00IFNdkDy1nTU8x0gH+uzh1+UGxuX1yRUxLlr+2cnh5XN
HDfNS929f53092gaw6PcJ8EB7W8hDZDL3y8dg9BlKcsuF93OM6MNh3rWGG4o180n
KJUhcaNbcjxJdPzcdHGWSS+0p+QO5iCWHRk56qhv8c17nyW32w93+URnBmdHGjR2
LkF6nj0aBTO1XKungmRJjFBWycOj5/9CMOp6n5M4yBopTcZTM53YFMFo+QQniv1b
ab9+Z7ejsWI9Ryv82Vq+ypwJijYn+z3q84AmZ046ZxzhquD9WynXSSJoQqZN78s/
MgAlTsGvAljQCHM6VdJus0C+Dp9MpM3SMOMbIqo3FLOU2lz2yGdVuCO2eCnOkvJ1
BRyTzwkW4YrZyO3QwJnV7HUkrgKr/y5VaN5DmT1aheJxRtVoUNcXz0x2KpdOWjK8
cTA/d9eqbB2iVsglP58oIzB0uznyIBMoo324vAeKRYQL/PACHeu3o5+Xei13iaNa
6C5UjiW7JRfldfLH6voH+TFOct4Xru1fbpDPuSW5DRzVoxW6etcM8mZam8qrTDS/
tbCkBa7fQznW+91AP3CJMmQgqDri+wbwG7/3yttUSjHHZyZCbtTbetNS8fgwTNjn
SC2aTVYrAWUycZMGVY0n1xrYr9ZzzGEZTX+7IZ6x5GX4B3a8LxE2zoG2uVf+Itbf
lsxb6nM8K+J9iEbOau98fq28DhSNOJRwX3GhclDPZeGRRNIOJD7C1jGazVLSOIPc
qEO8hR24wW5LTw31TGLWiRgaFMFhSM00E0g9DUqq9LJHc+M3rKDt/oBIiXu1l4ks
7f35XqDxLIlXkGMld3BMkjSs5q9KGvi0i5Rh2teAXqk/MkcfeYI9GdX5WJwncUwk
U0IryG0CUGHO7QUpHsqgUvluVUqXJhjmbzDyJuenxyBmBQ3XcMYPqmz+ib3Sd3LF
6hyxuXApj8ky5K9lDeLDWjYzAUyLfxC10lSjy5baEsjmOAw6KdQWTe1w0kCv+x9f
kNXCXHNTrCxMfcdLxqiZ6hYmGKMgKDAGUCQmwyIpGYSu+FJjBA1goP3cTNejkzWv
KVJbuGXKvkyn8vrzoLByRqlEVFPW2Dg48sYzloRZtQZOAEPWDVTJVvW6+VnpVQJW
c4vXXK18ldnstnO5EZgvyYwhqNikQkbtsATw97lzAlbQ5Lk94pmJQdjFkhGZ4QlR
fq1G6aWTc+3ETPzriS1ttjUrneDJZBYWai6scVCmlQipeY138pG5I+xmlOPJKobL
7ifVFD80O17iV59Pxzm72C02YozkpRa5UB2GAPN8KSTE813x/rEQoR7pxSwO4RnT
vYYO3rLmg+BI7G+/6t+4i6gJlTChf6ee6OxlJhSj4uFD1mRkgZU5XuzEMh/4E4zF
ZfoPTQsX23bnnqrOHBZ8EHB4VeygTWY/ic6O31HkV8A68Z7rbo6zRrCUorm3bbou
9yEW+IjFmJCqFIRjryLza0i+C5PzMhhEgaNde7wzA7OXER9jQ19QNh3QzvbqF31D
u778qdaJmkPc77VL9mW2lOuTMyvhlvWf/KkircgcfNoR6427tIdgHatD00YfhaK/
YHsFvsxrnZv++n2i17NIUkkBFWkR6X9oZ+nLfrwDkDe/vMpHnwHJjdqDIGRhvk8L
zaoSu6R5eiTDXQzuq6tLbef7yFsX0GiPI04OoFTHLSC+ZwI7uE2Wpw8G+avC+Wyz
ut9KFunWC8W3pMKrR5zpDz/Diu5S57J4d/JsM74Cb5BRG1RZXwIZSqNXyF1ekQP2
Ezdwtro26CvjWf+s6VXXpVNwIpjRiH4EGJHIeWhk/awctWtU7YePGHxJcQJPMGwU
PqOLJI6BLy7MLVx7M3piSR/T//wfTKZe7ikPnc1GcPGAmI65mOrLqAJ12x5bto9P
kyrF2VeZ5rvnEx5iek6ZgOi6Pn3UZCUP5PDDGldCWagEhetHO4p7AcknPqwPEcjs
c63t1e/N7zVgI1oTNjagkyN/sVfmlUbjPj+38DGyPrekCsTovyFUv1XN/Ek5OxU4
+QRXN9394Zp2LCLQYFPzZVqFchHbOcw/smYmSB3I4/v0SitCrP65tJU5iRnwPoqk
64NV/w7ga2S3eUcP36p0XdTBTsHnxwqnowgWT3GFrqOBoIAc/XsMwsq5YQGgb9m9
GqiUxh9qhm6eTWUrOxpP2rGT+gwSz+WlfYw9Q+AkoBgChiDzxDH3I6nWIPOWmIUF
CH0KsVqLeVSF76diGjMv/ynWTS/5aDmh9fVi6XPmPBSaAjTnrgFwL9so4KqO5JIb
xDPHj6ZRZ8UaS8A5Zf1kUzK+brA5gUWolnoto10L6btPgmj9sgdfKLxPTMTDxrTi
FfY7CDppdbXxobxLlqzGqnMa+ptXIaf2UcKXjc3q2/ccNkcfA6i8VorsTGgKT9aM
pRa5x65oJGPNdpdTGn2kNWwFtmal9q6dZiGApm91bGMKJWj3otmo/KWLAdj+KthL
+IM+PvzM4QTkWK6WiTkLOgzphQ+IWTmWxjVYYJ5s3SSyfVOY3gOvOw5u8hXpCzI4
Yy14h/snxd2OhBMTduPo1KAZ67BYNDUGgC73+ATuOAK39uAbbCDgSwa0eUqHjNHn
OGCYG+W0gy4VCoRDOG4wUqKIptPwuspyM+CEEDdD3l0yIF9vEg9jxbXI1ki8L9Rt
InIhEnsaZC9PLJrV0rf0Sz+e/t7ufAdVX0N2TG3IPb+JNT3h7vmUbvtSmcWb3dpi
HaP1pvxqPyS75I5gIeaY7+xNPFEPUJO7XkJNkM8q81YTjS2JAxsB+hG9m4EIJ1Ix
iZOFOH9Uv7z43TDRba50b1RFhJmXUGAlUjXogXrvhr8zCCJVZ6pHrTTABaT3Y4+K
EUryilsh9afZYDgDhNct00aW0j4bSy4voXuZZixA0CxDhBz6i11ojkjvJIqgGkhw
y0lC8TSiPFSBSpSgNkaFNysuAyE1Xhm7R0AnS7Uv1uVuTbeWQYGtDfSr2ADC/ban
kJx/x9wKG75xQTCgLAaUQwIa8lXrpDo+Z3RCAqe9dtsku4n23UsyvPWgifUiKkER
A3jKCZX9qQO+21Z4EcIwpl99bxkZej0mnpHDKq10VsAUocyqxNyaUTiGjmLA7fqb
02/fNr5WQfK8Y0DYNbDzIBdUW+gCFQd4rodDceX6wpzglrC58TnGaQT71TuR0GeY
yaUMPskLZbuBGy3B0e3tLUzs3nY1aBCPeFNjDt1OF5oJlpfjj12SpabXn4/CmlPL
JuhnS/VJndQN2UYhHfh9lPhfWKb4XSlBwFJmg15a6zOXOeUgN0QM+AvBYO6Gf6tu
j6BcnEXf3H37wJTS5F6ULh7y/smPAanVLzUqGD5D9BgLvK5PB4Q40Pe8s489Bl3E
k6UtOngEfLsYC5+0aoTNJUoMVh6aB/AVwk2HAMHGc6Vwr/CXCCCtVTrRbiZoB4Wx
YsTkx7Rx/1A4iQr8POdJHOS818hnl9JOLGm0hv68EMseMTgbbNfMd722SFEWkM/9
Dsixqs3WbhzsbqDd5qpZeA2LvhQFGOdz/sVUH0SJlrNISyK+uMa+VvnC/3WLCZRY
KCKlYCZkzqwlX83M4Szj76b8iFaJqmVSP2BpiOdmRCfteulk+kHywbWFj42Q4zxi
Q/B1LiYcD2ujdrVdkYo4lsri6H4G/XNPcH24MTXYC+IEq5UyXDARqbzPrD7f2Zkg
fmyW9Ih1+wqbatLZ8esMQNraIcSKyhXVqzPGx2dz9ExXO5gxaOFzmloMFMwyBzGD
aPxxa/o07zxV+7YvA+N6f1c+zN8Aryud/FuSvRBZgNyvthYh3Ar9zgcv/mpCXqov
X36WjwZ3KxZ+/gEqrJvsbth5gBv6go/7LoXSHoK0YuqkOzN0SIyBAM/bA35wpFjO
hiJnAR50oLJHEUoYpW09ZuU30nWEJlC+CQFhBpK5FqFOOpVAqAC/m4Kq7EwIKUT/
NAvF1ynoNtF8tEsXGjBGPHAyL6sxX4Nh+dq9Q79+03cO/qBfLeoi5zdwYR3uslIR
+mUOpEKU6nB18VTLlTXyS1nKGe8LHgL6OtRKD5KPWNnW0qlW/OQEKcwWYXwclp2Z
hIdPvlg2OuHtwFZoCWpLpJOcvrhDhtMY5Y/LweJ1tHrulFda/w0LZaYiV3K9h89I
5DMr/Z8G6YtnGKHWWbG0Y5Oc3SfxfNdVDRdLsvpYdy8wsHd7MZrIK7QrWD47JJio
LmZd9jTjj81j8T/5EAiI4nGFh7JCJCyOMOJceOe6seeVI1vO2OoEXPP2x2qqN/3h
ZuRLoYeQkg65BbNIJ7OPXCPWhNDDaFSvoX9SLAe0bIe1dPDjArpISF4FCTVFNEJj
CC5erp5/kb+kOVLlkf9LFVqqGrdzjBwXB4Y2YfSc2g6+2GSUZblTVzke7vauD/Yd
U8UHWugNVZ227AFYgWU3j1eaNlkNilJqMDxiriZ9MK0+4yzKU3NTLa9jW6wEiC+W
A8UW/+qK772EbAiK7Wd+bhCDOKF4Ym3dpddh1zx7CYf1oYXTIlvUZFJIdNUTJEyr
3r3i2F6adi8CPdY1Z5otNduOv2SZOwS2cDG6Mq29AVYzA3J2Qx7U7H/bbw2463Zw
6sAWv7SIUcbtpJUNs165WkmuR7/hrzVn6NB5BRELw7UG6z7LNYNILTMfG0hIWmxl
VRCIfkGJol872Wj+jzkujI4th0KBVYstmQ9CJDWIL46YwySMUS+vCRsd7GIoD6Ow
2ya4zoTLJxOvi2bqmAi1OU4ja5Vcu1LMejitPashDFsaRhUySORnB8t3BGQcfNtx
e6Dshzt4q91EKcBy2IWPZuRkscA32R8s9jY5sof+AO+9Dsz4Pddc6duVHeQ6r2PC
LSmjZbMUTBASdirJ3bjMF5P2jySKCpye+Iy+xorQLDq8f9huHrpl/lYXO8CiBNgk
lRXaoBi+zKuMmK7stvvZIz2piMcUnG/ET0C8ZjYBz5gieYNs0EmbOI3QKpbzUOAy
pgfy9qeuBslnRfelOJKL5DaF5lQMKgFxKOaW478rBkExoG9gfbWKf97CB+Qc0c9N
QwXtfI0jM8DT/v3swgwJrqSWmg8DnPoZzzfSYSw8PKezg8RDjv3FYz4/0WEeBcjj
fJeiwBQqKv1C4EiUQbETKheFIwkLPTEJHaPFNjjamkeYpO+RMQbyU0vZJcfcFm0q
J239g5cQWxVNsc+FdQnVrtE8FeMIsvo2af+oBIwOjgXkEU8iEGItbujCKaxbplXQ
xRCw02kz+bl8dLbVYDR24BW1OIyB+PnH5nc/JuKd6Nn7aNezheGL3+yJUGZcLR8N
aaVv5gt8s149b74JxdUQpjiTKt2O9oDVYClV7buwb7eLO6Pf1kbFKluIcGKH19oU
JIz1eF4AGWm0eKVbNtICWiMjUQ9PSRZf88s2GJEPN4zVmJEmcwBF6gOiQPwtv75U
JwaqQCRKdcBRqb18j5gs3LpNHhfF3Cjif24KoJcNpnXpO5/pgs9Dea4728pAcqDJ
FyQvJKuCEO7U2Jdagwg8wQiPyr8Frkk43pokhFZq5AYpAjX15TZJGatclJ2ViyFI
FvQPUyKCLHW7A4pI1hAr5DpSXcZC1FvIh7lDj+4et1VJUjurd5H5IFSsv86emqWV
+fiNxuwyuFCRJCF6o29aWaejgxCRmlBt25muPrfLTsQpSlCtXtS4YzyB6PuOTMy0
U6z1F47DiAXYo/2qBlZo91uC1moV5akyDxNsQiKZgrCVbn3dkthoVrImn21o6ZTQ
jxDNPO+Uv2vOj/MOeGETW5AMTergeF52bc1sxL7v2fZAsXw/Rs/zaGUY0YZux00+
g8DI7Ys73dP4Qhxzlj++lsANUvAuusoXY2JSP0UUbEVB+xZsYR9iBOU9AcDzwUzw
7fVWi03f9phuKHAKhDoiGjhRtduUbuftuzOhLWVujf+ktNKyLdJdQ9vK0W3q97vR
5GAvItXLbxap/UZPx1+srbD4feJWRWSH1KyxOgK4sRVn9gE8B8ebyh1zsILSSdA6
I9p3wZepfDZBxmK9F+Q4RY5ElWATiozhBstgi8HRRwCNRLHmfX28CWUuk3aDnt0n
mou74LG86ra+3ZMzvgLu4hniBdm3DSUtnlFF0vqjSKRDZmfY65u2avsWKvjscRCR
G7oHEgUhpDuENNSPzveEfWCiO1sRnleWwpuxXEfSgsCX5PPVkoLsQ6qKE9Igb5nH
acWrmmaK8Xe+8Wbo/G8LN/qtE2sHMpenCJ35a/FL+LXXsMVEoK7q7GwiP8zfEphy
uUiRaujL2aKLhHY0tSaPuCbE87fNEGGAfulln2mflSc4virz3KQG1zHW+vr0mEJN
/x39Y4VuWjyYU0eldu2/pMYElvty44aZv67OV5F2u5tbvYoHpN5iDvrWB+VgQdUv
vEfPMYMKmCjeQ+oEAKYSg0rMr9AtJjYj4TxjgSwkNs37Xd6UHtjS1UndD7EuxFh0
h2g6L51onbXVd5NJ0fo3rRVEjV5o+rIjg9yxCT+KeHMnOSBeez4g28rBfZz4L7ub
oedBFMxSdHS7q1kHkMGIRO6rNoyAMAwRzxQRY5DfrTZ+G515S5Y07AvyWTn3dK4u
+jx+kHLk4RRptaJvyxqP/uiPJ4BhnQ/8i0UcYwke1ofjcHxzc11iR8NhJEW4kOcD
gcg8XCMyniv31E1EldHZMnmzFFrx/DN5slBJV1Cme682+nrDx9uC5Rd+4yZK4V/t
kghsp/EeX2gXYzFd6oRmN/pj66ijkHlYCFi32DvkU2C135Afd77LvAF4Fh2VKM5c
Pi1g84++mkgjX4PYg2K6qiw+pZ8MgKYbdB5U6DAbhL6XlW9dd82L92x9JNE0JqBl
NkxXEMDhVz1ejzPRlaolsKWPGNjls3BF9z7Npetajnhumddah4rQfjAJbRKR7K/5
FLvTkPX0EjQwGk3dsGZxdWR/k1tRP0BK4MHwiHMexIlVhToGRnm3T1ZN0V1qfQxT
UWXzpAf2sefADZPZpTa+Iv3kAlH1klcyrma2Z6uZ/LyyzOxmFWn4yri1IUCe3Lbk
dhDKmF9Tska2r+tZta+mrttRtWmG4jm1CptbTCMDKtWeECJXhjfttR/hZXUTp1LQ
d9qizxZYkl3NhUzXuXn0FQINllpJEvbV3U2ZiW0c1QZAKxB+bjb49v+lXJ+sru+6
paMnJWbIkeHPtloUbH7SWEHflWKJHBQEa3EMib8L/i3U9B+tF9/NBzlhjjY/cRZ8
Fky0IKX3MT04IFeT2/3Ym1BTvukEBXmB6ohyAacv0e/iN73eulIjVMTzs99tnlgG
tbx6aV83XLrquGREQCE7SWZwhG7UEn8Agw2HkXMc19MllhuXEWQ0QD2OUwgL974y
2X9NJiR/4nmDFkdwz7j96Zm+iyVQfmad5YL8q1qoc5nUhAFAgroF21JWPwurmkWn
09/8qq4e9elIGiaiDvVp03MooqsAQBny8XDi9YCKP79TS7foQYpRtSHXco3Uz+MJ
u5OTAptdXdrxV2LHfYf8WR9LuKnIW5xrhz5YziPCU+XhjgasnZV2FhNBRvEeP+eN
ElBdMNjaKAw79vaSB1ZSh1ZnOv0OSCYyzFGlKeXdLpB+l4pSYa/R18tmbqorxWwE
Mdxn4SsalaXGQUsZqtpILEzey5BeYwXJZatCm2Mmu7ww76CZKu1lfuirD0SIujYB
Z0XVMAT+jdSDltQ+NMeYqWROo8i7lCnX2B3q0yYNu3t0EV5KCcR/j/1lMoYqL7kI
XZyF4GmguiTBHAfCJF45j+lZNWR4mq+2gOPYpolS3kzh/ULk96+isxmbiouJwslT
3y3NiYoGr21j0itOOTso65p3pYx5K6YodrRz6PyVPkQkvBKutDYzLwbraCUR/J6v
ZhY7dU4zqcfBqNWUiwVw4RjrGl+AlDIcWuVJJ16VzaYwqSFmv5CBaVESiPCcqLih
oQtmkRkHRJT38m1vqlG+Cdy7VIZ01Enh3Q5oHEbr27p+OrUVnjcf4QBKpjWzau5r
ErbeTv794tER72LNkb0mppHhP2fddHJjOS0nShMRg9sPWRGZigk4BZlFAoKVFYQG
2UeQPj+4o8DrLcSEinxDAryR9EUY4ptE8zGIBzDdQ7lHYHoZPKrDT2fIuD8mRugD
rTC89ZQQh9CPvaI2TbJtuiAeUkH7Y/B5vvk0DCcqeI0bZoWJEYVTSAEHnYDaM6gz
2nTSiTNpVuoQnz9MS30RtZ9ImE8LMyl/87NpWUclR3tIoetPsnrBM8N57DvsiaAS
kUfq9dlw48vO0yG2re1jedpl1QYr1kUlSQ+cf0KRtoL/XxZQhQuqIf78xeH+QoNU
STs6z4qKbw44YYl1csfqesFLLtAnmJ+6gXug3KBrInRbhBgxNfbh39fj7LQWga9x
WLqoiOcdsQoTauM7NqzJURphFPY5cZheMafYk/q/P77ZiliKWjPFui3vSTQIAUdF
WbBSYno4j6YJkR6AvsOLK1IfGJ6qvL6jvbNWMycIEcRbw+Y4cGL4Tf4ubGbeElrS
IAREpJWge7BY4MVwFXiYiE7hfaz7gBIY9e2OA6i7Fv7RKanavBS9ED/PMg0AeNCW
QWbT3UhEVvEk/ns72PKOCY0SPwfOSUESFjjc8F6819LI2GoZ38YL5a9VnHGCMI+R
fOuvhY/rsW6Qbqw0QXUMz886yLdhADBCWZ/out1nXFQTXwzE7mbg1NVPL60/QBeA
ZZ1Q+rY30jbSXHGyBDrlSNcnRT1yID7WzDALfKjZuyLv0Axt4XAzKVk2mrlvXO1V
DLlwQkY5oaoF8ow1vZ5hANZY4mg0qkbU/Bssa/ESp1UwwmTAAy7YsoJwXnT5Lu6w
CVU99W3+lbqXtUvQVMuX2K3zr36QJC8qwt43rUw93s6W4zvgjxhDRvmh+b4DxcWS
wfky6JyTmefxwzrf11Lcp2vE4fubYWP93fcC6SRGnF14iu6FKjYAk/cKCYlxz4+B
zjolQeCFDSbaNnU1Y4Vc46qWisaUJu/cI36ewY1pOApHJTBc15TUvedDX65nAIFi
u1CqfRQVgNHbq6BB8gDhVfHzfa8nPXjlxqaMKESNklKD05ENLm/bEfWps9C5u06X
wbOl600qXYzzS2Asy249uJlOhQqEcCoBuGM1rMOFy8gOEGmlX+XMZrb2XXvV19bG
W+XBCWA17yvOWXEt98Bfhj/rMZxSqaWdshRnx760BYA+hpEnqfGgC62gwD7lR0pc
BMgZ3ZUXR6jei/q4b1nltFD5iWCuPjNgXzraNVD2HrHd/Y8NglLILF7pP5uYOl8p
qTCEYIcVVPKt9YziPUq75MuMwS7SeXaoJTUSwRnVGf24ZrqmeQkbNLIjXS/PEUdH
Q2I6Ec0XfMT8trjUNWHT65pGm0EW6RZSau9TO3HTWZLG2z9BHJSNJhZUKeMs9vQC
9dcHrn0yZ51j/Tn20Ar54Zdv5UjlpCbQ9LL0kXtoRfWt2rE6dHhA5tGoqhlVuLpV
hYaOHmmsZFiXSpjKF7IUxoYDQ7l7yIEknRNAXT33AGUiwk1Xu+htgo/EKgoWKkct
aI/u3cVSvqNT4JxnF1Ex8YUYWCyF5iXnSd1a2w/voMGQOQea03+Hhi+omAzhs2xy
GVTf5I9imJk15WBNMDmIrzAMWH8ILBbiL/Co+3TXc9pJDjjJUandOa4iaQ/slGXZ
Rm4S/gmY4MCTWkBYl1gm65leLLl56J805Ws6Rra3TlPoH23StmqRkGcx5ZymdIaz
W8ekyQvqnaICzMSeT/cudlRNEzBsEnzZhGc/vdLhO2/XCj1PHcxfNLVo7QGrITkM
JS8UrrvEfjdVW45yhqxU/z+2SINUioohagu4cUhDSYN5jlt5Ug93PDn45brluILo
nCn4lKez8qjwIrw4IYKdSTLzOUidGbvKMODmPmricLN6pNoWhrsSf09IcKWalv55
yC17bGLiDSrkhWYkvJGvaVZw7eKvTUkPHibTJJB6xspUF0rEZUsXEm12bkszYBTe
JpH5HHm6a8VZxZ5zWwyFchxkn3J9ySkv29NIUhblh27UK526T0QOfKj1TVH7gBwG
aeLMn2kUdxI0upRWmp0qDGoOBxD9MWJWVfurqRmcCdHn/wbRWCcpCJF2ZQBMKIag
zmow/CT3I7dkbk8sU1mHtQoBK2FsoR3cPnx7HPfPY6lVeulL1JZ+82J64BDlGyYh
vd5J3KeQ2eJt3I8vgYN5sd7S2MpFeKRpq3EIkbIxPAEW4Nzxn6LAdsvFEHXtDlBc
g0ljFkh13MPFYpHra5SnuY2uogyk0MG9TAKeF4DWsyeRFfY7de4+5jflCtec9e40
Ft/nulyqtXs3Toh3HPD2ycHQFp9MyGgFvMInx+rWVXgFlP8k/86ox+xbih24N7bu
6pwcHuD4kabThkYm++BoUzPLbf5ma//S2VAiBcCTS7AboXD1A6aKsVJqX54oX0OA
0Iv3CFPflckbPLbnQX4qEMOb62wwJByh/3BzDayXFvfNe7CRrzL0Xm7sqqSqCZ7f
/mHMiA7/qVKjvrpCuU4ok14Ovi6lRQJQqOs/CXJ/RqP6TKUsQ3h5HHrTHn1SLB6c
YnVfmK1PeQoYEO9ZPuEBw+gKs68QPQTjGenWHREYnyiJgv7n8XkemjlKEqWtM3Zt
wyqKS8V+ktP+slt3M+oYA9RUCHjQplfzvCSSTR7Rps22z2Yq+TDQGlrzuaGHRegY
ZzRDoWTKAyCjvB3mFbDkgBSFmY0SXYGU3pMlrgXBp4C5E7zrl0t47uAcpCt8Q5Ae
199CL9BUxEMez8PARud73rkSnM9z19ZPMUAnBz0az7OTiw4aIlXdndzkHk7i/JpN
pUv0+Uo5UVyCi1UOwzj6FcOUqFeFXO+VKcMVRUBR4vEKbAfVPT0EYYbwYeQb8dNO
XbeKF54z9TqURuuC2k/hzy43sePnPk+hXZZ8360USr0WgZb9Wk6EtQ6BJykiNVES
UNGd7MEH2DPJyNcAxKqT54akNbmLBhDUCQR2pW15YS/1Zz90/e5cBrRB9O9BXpRU
tj1xgklUIjuESdysJq0jkb7FN9FoGItMjLk+7FIkT56e2qt4YYMkatlkb79Tm8Y0
X/YPE8Thq/OWlvmxBzcqxc0pXge96KW/c+iLJz+p1m5ApNBBNu6qZv1vg5BgLG5g
u7aNW8FkTjrHoY5tmtnlmvUiSg/id0zaYMqHSyQm1XEOHUsQ8JlURiNwpCL0r/wv
4gvSSgsrRJfm5Dtc/KPx5yxbOuTRVfK135AAAYS+KVx+HzGHcaAAoRde+Fc4DmkE
4lhJa8qrn+9OSaTUp4ioUg17sGt9GDzsDhoWk73XTKvYdBnowfBR1ldv0SZXkV/f
GwIH52g+sdtusDQaev1MbujBrpI1fs6J1No5hIK+S6BblBXevvTKZrZiJjtHFg50
AoyT8698GRMpoNcA4lqmd9qFkXRR7uHD4zE2selDYZExqQaNdpJx3BzUeif8XiVg
NBfNQFOVtcOLcUPcL5xcWUoFOVy2zXxh4104Twgq13QoOWD9/FnzWYFJhJ74nKOW
a6I2Gf3lkMaGTkbfAs7+GzJY0FnLMMO4QHF4fCca73whMtkPm9wi1TzybLsKYtMH
yO+mYW5WxSZH22h4zPtHwgnKgN+c6DG+7zqmDnUrPoH5oJLyQ0GcEYwLcH32ekle
86wqvO9mkpJQ+AxiOwdagWCRbzg6noaxNxL3yljBcUaiLiRWGunP7Ejsm3Dj5cp+
egDkWXRQe/AyE/IfUmmIo1DETii1g4GoIyy/abAJZEqmfLSVfn56AxWvuJ75bG5v
5fj1MLl/F660PWYpT3i3GxivFHV+mflzvHLNxRjeqOeCskxZJv1fMwyRovOA99E2
/W6/6O6PfBiqr07vdxQSzJmkLaVLUncuIpoy4/lr4aqQ3T3Rs3ttb317fFCGmjaB
ggr3tW5czIaPmaQorFX0wg8uZxDe34yz1EeAYjjxL8WHtLcvFQ1NqLDwhzrpDj5w
V2avEF2oMusA5atRT6FTfOGRiOPhzk3zXuLlJHhEweCrUm0HAMxjLL1EwHm0oD5D
LV9uNfX+XlcSooJ6VHGCQUBr2b8PGLfs0I5FS4wbryhV4fKLLTtPltfqmEgCJvmi
DFL9K1VVvDdrygv98xdDNXvKWCn8Q34zOj8O7tOzjYhwr2Z6RTBjAoGOGbbZo/rx
hDCo2MhzccD8/hFrni1hjNQ2KFrBW0PuqecqlzbGu/wIjtmUaIiOJQd3rIzmqywE
L7gM0iQIhZzZ9yOorOjMLhTQgGqbXtXTtlTY+IfnP5SVg7N5FL9y/Zaenn8Eh5bA
EXRZKEswZTjcy/OglWzY88jPf8F1dbA0tna3CjrWrPwiME+KKJOZ+0FGQomLo1bH
ZvVbZg6UmWx2q9bVZV6z1uROU6BFqIIGQncDWJ8eK7lQFeXaD2JMeug7S6aXZmBT
mj9SYz4AH3k9uGFVi6yajR1WV9q97pf2CwerzJkwycSUj2JPHVuGq55jv6znYIzo
4y2SomaDA2sqcLCWGB7tneqwftfq9qOyqDTgrW8olak32ZFn9pzEvo255rI3ndZ7
DyUyIaNskZMBWjHYovzXSjUQ/Lh++2iR4SGKfn3AZEN+NVU1opccw6Hj0xKwFuyK
J46Z9egq4T7VJiqKy7i+0yScF2oMjQpf5DjpyL9wDKxmf5l+xU7e4sNeZkWCnSM9
1yklmclBjO10uBIZRMTZ+GVgPV512YG2e5tYcg3bNwj0KGJygwt5ZIfb+kuGItV9
jOb2BdlWdHuYa94/QTPbABOmOtLyCKGCKA1EnW2bVMEXxHVEPbrIV2OPEYi0q6jR
FXx6GtFCVdcaAjDD2DCUm9a/L3u4JFGEFWG+eGfMi92Btb6PvNpoE65QiWx7QtDI
Kur+ntCbJpEPMgDSdLx0E/FNCJggFbSJHT8R9uXb5Z2vuLgbNGAohFR0S4tmVmhp
K1BcwWabVEtlD1Twp25aLPdGpdUHcSsuHlA8JvzAfBASDbSg0WXD/hOanka0nThq
k/r5PZp5eU94M69IwWLksrr4UsHF/U95txMlBneEcf0Zp7C40va7IyPCGl6unW8C
zJLE7/qdWEcy8YmWn5cW5wjXiNSgrbc2pp63IyFqW4GSFV8rWZvxk/mkQviy2j3n
c+ixmAQV/iwHCX56H4AcMvfB3eRici/drCtqlUxPMl7exSEZbOpcdHytzCWUlH0o
KLO2n4C6YNd5uis7Wp8stzgLhhqCK1Of82BNh/coMUYUPFZYXJ53PrT3o96ZBTbG
P21msdJmGKbTr1eP1P1i8wVYYlE8rjcYXR7OFI3XTzqh1rBMhCl7rb8W4tT9cA5t
IE7VgeaRySRnCDwhpTqqcwhSxVVhZDnrStztkgR70JZYzlBdryMDGfieL8w7PC1n
pUHQ8Z4eT10a62mBnVmFtL3n6VU6jbuLgHIJ8J6iQgvhfQlF255AkOadr+CLIhx0
uYelq5jU59yOXYl0Hlz79nxPXrWk09rxwS/hFCr0mikwhj8m1kUC2n2XuxCclL3G
83+RYMztFuivYv82KUypWrrFGwTvJahRAGjho6HLzja67BFMwhRLz+NEgw+W+vZf
XArOtDmliYPp4YUZCKceUHQm89z1T+uW1lA/sf46SRpupfOLAXjGJiyuQMvs7X0h
tnABJ2VyovfF6AQBJ9UNYU7M+o3z5ZgVAbDT7scy/r4j5ZyANQE1Bkb8dRI5uXHb
Qhe52dqgXznaUSEXeSJwBglE9HAO46vHCZtk/lIhCxZXFzMYvpGsVgKpO1jPztQQ
1TaFO1aXmyHQveq5L+TGXcv3+3bMh2enX2PdqqzodvqUp6zL3c/Bud7w0oiGNSZz
UCapAFO5p1haoemK2dZo9pc7NhlIbhXdMhIWO9OT7Nvp6zYgLG68kw7yypoFHmdW
spblPTGRULL6vX7l0B6S6plhtJT7ZAdEsBcdftPxNQ2/AR6dZjwLgnctNhEgiDve
de9mkqGeSoPIGkw83Pj4iPzcJiBF0dxaevksYHBpSTS4BSnr96Yj9XN7fVKqp3lm
PtwF1oVKew8WiD6FcuBvljlvUiviA5oXOSVFB4pITsQSM4L4NzsS+SVvCieleyIG
Zz24Zg8C+UREgrmdUbyzkncwPRn/w9rMx/yI/K724QTDWc+TWcwa0QVOsMvUOdaa
GkGBA/pMH9MEcLzHfza4TWScoZ2yy0xSn8G5DXaoGjQEdu3QJRQlXJzf22prlfGU
0OkjTcsTuIXBSUfLbNmMF2KM6S3Xbnu5m83FYYLhI5h+tK/XG9YE/2IPVaHL8Ltj
vhjnrm7fK7TCOorAzZz/crAWhqGf4X/Gw/IQWpe1UFVHZZRh44k3L7/LhEhxsYF0
W1kvi/THKK6LvhBRV3AdFWgk0LEDkYCQDz65/hCrtwmMBMrK13ojFepXQkHHVRjD
CWvHzwirqG/D0H56QsOodx5OKreDmkUiuKTRWXF/mq2Qh9ufX6n0+mPokmW3nJpm
Q0WPk44geRExf+Ppvg/lRXjNQRbzoecUnYa4jGXsh+JlZ90Zizf3d4qO+t6JCbaB
cHurJoycUe3An/aekf/7veDl6Y627oAwyaf7w6W3OA8rcvsS0Q4ScvkJD4womW62
ndVmzIHg2yJ958ctA1nvSl4dOTVhRHExyXQgXPFHKkAtmnQM0fNGSB8RSfCJguaf
hqb9c3sypipSBUZwiEdqokSE0jK4v9MPApNGrh/pvPECDqVcYmciwVIUYNEF8jLR
S+4I6SWvmEgVz3UQK8439iLIq8hF0L2E4BNhnOJjpJocOJQoLBRsDsRSbcpOoBIH
1L2tJdaFU7/TqJ41SzVVvZGgpZcBKnazQcvTi3wlH/J/pmVan0++bD4i2rH9hyQ2
8j/iwpWqo1fdMpEqmCz88Q==
`protect end_protected