`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 4320 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
YachDS4bpHRDzLXFQC4CtbmYvIKKgGLmslhnluyqiohCrDBedbYpvxvawouD5zIs
wDCsvebxutLGEyQ95hDszUMlb+6kepn3NMTpaKz1Ov3IoCGUckNXmfj+we0u3RGB
sBAhute/kgpQ822NDFmTvzLy8ZT/BMkRUXiKbD3o4GDRrHf8wKEpOc/BElWCnVvP
Qs+uXByWKbYOWE7fFJhUsn94pGBctJHQskoJz190GjiNVsRtji4dzcnQYJfIhadc
wbrriNJVgL2hJuQgaGlhJzLMd4QqHZ9i3K4s0k2hM3MRhNEjH+uo63jGk0CTtTTI
UkOX/fytroU79ZsjOicsRVFhwWUoFHACM3JwvSbKK1YzAkoIsF13IE5SCDKJC/Yt
ZSWspIz6JWy4dlUUuGjgRsoks2QJfMPoiOn2VQZed4vDPfXmdwfc8cnNol7mkeXF
c28QFadE0qh4A60WwWQZM5rDAvX0fWK/8dAH4CCFFk4OqmGnxen+KGWyTG+uNMeA
sXLVhiPVPqiNZpZWVzg8U5ozcx64GY3Z8lAOFcml5+aHGh9Md2wHcQkIxgw+cYTr
ne5oOhnnKfTkJ1JlzLdy75S/tb1p/s+FmEXgMEU5alzreodzi6cuBp25paWSAXXA
AiJRpmPW11igbLREZIauBYxNjvTLGn3DM2iG/NLMb4shbfuOPqyDdfUeS63dnqlz
CjKwOy4Sp/QBVGD23av0brIlGBGMaYpwQQkyEvblQKzoRnjsMR24xC6RkiVbZkJO
cD0FtI7TWr1+dFyOoo7Zc9iCqxg99i/oBiRnEAcM/BDt+MS4QKata6DrzOLp6Htj
bfLhCkI4m12eZrYG+G/v9cmLy0FnA6TNJFHg1IqNo7bYBDMcX7RRWEGciBuGJMmO
ISM4c56PIp1QI1mq5Clro1ADnE/SJWUtgiPsbOsUo1MdcclUzmGkM1sYOl9jWMLy
ub57SM4RYrrZmil7hRDIU+LUX+owoSp7tjT56a2GeJx8YKjgeapEYRM2Xv7N5nsu
RWubJ01sprSisJkcOpcVXw2pwERb54zi7ISH/ecNAWc4LEnomDbqYsW0IGy0s67S
pbBVTF40XVtKAFRX++I3ZY2znj/av1okDfD2lkY883V9fyrh+Vkwq56wDqI7A8VQ
qUCIDTAH65hvWAsiTgLFT0849s9DxOkdkMJIVe7tOz8e+zTKaY5ewBTduib097iC
2w3HkaXKhWnx6xt1QmyLLauzuqk9+JDBZyzuSmctmSxn2gdtPxQmbAw1bzR5jJVH
uNncogfBKmxK0kW/6NqoabEW2pu84wSTaeDVihRbElHKRWg6bjOMuR2KZDcgVKQ8
RooMpCQF7z6/sYXhgDCQ5vp5x8SyNU+TpotuwRX0SVBhzEwX5qoD1xa1NE8OaAIm
UdeGKdesN3mOj7Z2/l6qDXT8L8t2Ij52DJU/PFZqsmexDwC5qlno0zW1IUwSkozy
QGArjgRJGILroUfl3XL3l/WimdSPPJuL4ZY9d5UeXsbmawovgkL7bqIvePPO7YYv
oEHV2TD9rKfaq4bNHlcXpznfE9tECM1L5HDiSu1C9FdhQk3ZQ5EE2jrjCkFNPBLN
RvquhbEaovYXs0nhxN5fK0P/qdVKv4jo/Q7a5U9yiX62fL+to9fZLsRSQizsGdVn
l4IBDxPatcybKfPizt2fEIATq/WlzpGyKozAJR/looio9+IwcNxkegn1XSjJm1Xc
RydfIdXule6gVxct8Xy89u+lDJTiKu7OJjQF4yuUazOk/UbtONXlaNIrBgKyEPSb
fbJx2xEpezBuaAnkIwaIhgBMtBGDheSGnjrNkdMMjcuHAg9ABheS8C/51Tupbc4e
QRCZ9Q0NUtPyYv6VDO6keC95JKPBL5eLt2kfVKZaFt6yHV/S7EjEeR04ZCxDwQ4W
2IZYqweDoWXxprZJfwj2TiJgCXaczktdHTUYIHpmw8DAaLdW+QF8PfZGjQBgYzMv
Sw2Ox0od1xK+2+5IWrqbGNXBkLUtZSiEAg6F1Pf4E1XwsX0cbJVFn5PrCjvM9Xz1
BNTceuIxc1ymBjmo1d4fdRhELpCncWVSq8DqXkbhjGGxxj3zJP6q/tsWi3WymLrz
SGFbiQDT+89Lavb0fqSgpLTrJIgQctQ4+9IfQLo3V0mvRVB3qgyi+GTA9psNAVKX
plrzds4l76xP/cK2bUxUQGYD0VS8YseVO3bvPERIcjN7GmCwF2kxgJMILtueyCJC
AeEWINFmVXdRzDeuEYbI3mb6oEKXuBq+oJnd4bHKcrgPQXrrn4vgPhH4zvy6+oEP
z8Elc87jD4dsaqv0dO1pIodzOJUpsge5Xrrh4Bv8aLAwJFE8P97ILz3x5uar8Bee
rWcVsH+czj6eD8RKsWan7r3dy36wmJRk/p0WtBKdgspncQO2mZik3+XHT0M9+mQS
Ea85P3/l3F4bNK7MABLtjss9ABa3AkI19w82SXQLGobZ6AIExhupzYxQyvYStwhH
iGxzQ8ooLzgFalRF3yEvbeW1JrbqSQA/p1d3wHAfAKUWUUDVJrlrYFqBBwT7eZ/8
wB/mQMA+3q+ULhbdf2Uq4fMFnrNZtV3Kzziqvrz2jjTwT0rKd29iCw21wB7k49Z8
8YswhyzhotkEOQ6EXWJpcrXfMalyZeVo+76OtfggfzUcMQRCmgeSIOpmn2fC+E2+
zsoXeuwOlLI6aVQ4q3YWfnXDP7+frR0YNLgzOzlRVps+kabPzz70nWDHYa/7pgBY
IsGFLWNa4MXKkVHOyRD4Qey63H8GX88yVXRnfKuV2HZmp2idTT5qkk/AE37NAxOB
p0ai6SIivc4jHrsU+plsNcMxTUKsfkTgqUXg5Cx6qfYZgwGOnUYa6ltKUJi7f6C+
IOHQBWjzlyQXniJdm2NpMfCbPqMAg6DrspHWTZZhfBMYr8ln1vn6yzWz98wTsCwj
dn3PDEtVx58HA12k7ESeZrB4/BlMIfM+/wOtcK7erMG4YPONGpPIAJHXwGhX2Hvq
v/D419SYbu9K2URKMAjLAuwOfadEt2qDXgEBD+bwLCPcYz9mzjbcJp/54VFFdO2P
paVkHJPkTJPHI2QaosFoOrxqTiGFBpotqblQ/qncU8b3HbT0iapXLLjPHSy/1DQE
oIBwMmrTciXciFX0GQM4otXfkUKJdIHsl/EyEjHCits2SwVuTaV/nXyhUE+dE6fo
N1+2e2qW4ppI4idUZH64Kfa/7EhXVEQBWQ3qYI4qJh3Yh8keDRxRdfFLOJss86CD
rOFwTmoc2PZX1QUH6QpACj7zuoBvzbi1lSL7uaEe4Sjek6CbbAjyhXIJj5kXvh2K
zpbkmqPM5oR+Riqj3CrDOM76G5ToWDWOG09g9ykBXlAGPCAu5uiVnk7gYcU28JMn
FwuYa7OYEXtbqb5NmAod9ycbt7wdmIwPwGRn+3PWRBTNBMFWXYx8BJ1ZMetoYWgx
nVtBqvY2fp6Mu1aFhIVXbEKDHcMP4U86y7Z3e3CLwbQc7CIE+bPQ/wjpU7RUNv9b
xUCmZTUWELXUodwHyZ+DtM+3fxnRcG3gkfqXKKB8KpVtwxXyF55lc3pv0HERiPnA
8BWY8Vsjo9Wi+Jju0mcvOvQftvHjGCaIqzhPAI3KPQ2X2MA985jZZhA7Sg2XEhG/
8e+egWiY6cdiE8LRfJ7lw9B65jTQ1U7NRo/IEfpVIYm5ApQ/rdUhmdo5E5ELo852
sNJf9wjyplMjOEE6WCjtKFRQA05yO+UEN9g8sgIIvYxe5Ei/cWAaX17pgFKP0skX
NDCXOOeD7GB1t96mimxxypHd5IedUR1itRCqCWDcpVCM3OvZeQmQGPIuzENXK3WY
OaavGGUDZ2nDl2D0STIxpwcCXSVLl5H6fyaoh1d4FOzpF3s3gxL/jregrGN/PEfl
wMrnxi2R0mIIU/Vq60TO+H099AuG+uaborMvfuewuds8wyDJQWvr1+NJ8yrBFt6S
BzjvDvvWYur3vgKGM45kBGqsiVh1qUWIHsJFOUSrF8WwfsgZPnbUvFTT3jIiG143
BKi/+B3SC0keGoNcedVbABdMdoEQScP8LxpeeVudHJgv750t4e9DklORib2wyFgG
iGszctZWAwHuGZvWI174+BJyej2IRcgnEpUQiz/deVCUxeJulygSAVKXL3r+MULC
kHdlQiMBxHH68yF7mKSTSWHtIroHk7flhaKMm3hSKBZA+hApLalJDbX50tc777Io
B5yqMtkU3ICCVVbqYKZIgQsKa4nNtZN6UGmKmxgslS2ukDQV7oCyyVGPTVj1RsZa
NXHjQhB/e8i7whRhpTBDleEJ6HwByHGrOzhKTVcO9fSWRyoqiySM25h/WEga59k/
mYV+0mhWeP7ccR59/n9qZGJm2yq43FwqgKyuJlUCwlxedO5M7LKP8krTpZUkD+WY
vW0d8OUi4SElmX3keMRY3OCwzE3NFe+PXk/aZ8kIb7e5uP716Zgp7iQjaodWQxy2
RiUtDvcmecEXadqVa35KzJbG1CKMVf79HGiPPQyOOp+TazfSmg0wbB9szhpOq3W1
4IojRWZ+stc7F2DFBy0vEmMN0/TMFoWPvgQqSLsfK9etm2pAFPsMLmfBA7bn8hHG
l/fAVx88uh+sck0nfN38jXEvndTDyJqLX7+OA1ovVQUj3jAOtYvHY3PGjqoKFA34
oq10CJJ/gcIrrsKF4T6x1kzjclo8J0NH+WmPILgNrldrMDRn5+QzSv2aDMeme6ju
UWhsar3hRqTaCk+GyKdqJO/esszSAeW2B5f5cr5AXgIAVmTWNqQsx5UYHgoXyqVl
uq5mblEmvgpGfNlaKlyfabyFwCk3C6t4lACmfs2Nv4/Lwt5T+/5WQqdGs7y2BKDb
D+PM9wMbs54+E1rVV2NtryuzOhVLiwIXvyqyjWMIg9c+qCwXWaWDhRfr7/BJHnXG
8p/PrfAaOUZVsOJPs7359DrWwrYxeA/E+9g49SCf1Sal5UItbOicQuIa/yk3/oru
8Oa2hH2SeXpKMcfrFAjZPJob9FArCwXK36Qdp3z9RYVK/T6OVPe2irvh+iQBCp0H
MPx704+zFX8TZ6aTRhavaBJEhDCIftur1rUGtiZMDSUA6oN4fKIvSZrppbXyhxpj
vloW5l7fF2LnSDvxeiEojYVsGl35kXD0bJ8RH/ECSsHBK3F/jjbALJvuW03UYYr2
+MSL2l2RIndr2Hzc22tHQlLQpml4ca3egsWqc1GrPjTiBzFGx4LOMAlN6qixA/5+
HpjlxLxowsUQSOowz8F0Y/ZNmcFOEsSMer+9O7C5KAIVuKq82Mh0t3gZfhD5Vj9b
l7U23XnAC+ivF4ori6Lc/Bj7mQv5mICDaz2DcRbHWe4z7WDl0NbwmYopF49Qa/xA
C4Tc7MVYFYvqsFtF3bKwh+oILghlsjwAKiwCDgjq5GvwXGoovNmT6lz+Er2YkYir
4lB+cU6vhYhYq56r4i8P3/7T0T9DzNajIPHwJoGmKYLHpSStApcMvVW4r36Yhoju
qkfD53X7YR1j6J2FuubObtd51yuLdybYzRsJ7IPPwRgyLg00+yCy4/9d4yQYjw9j
MHlqDPqoyMUQQVHsucCjOBX8WH+oYZj/TpYo7FTdN6dX7EEiqCwMxlWpCp5OEo3Y
`protect end_protected