`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 23952 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
S993bpJjwxtMDn0RNN54X1MSvtEYYT/sbwehd3VbjB9Cm8+xOsXs95knYAAllqYu
Ts79qaHImFtFaCU2t1vTsaUZ24Oam8qBiy8WKy1pehTmPf/vSrCTygXC622jIeiP
vSG0LIna6QLXJzSVZ5jkQHkzrpmfjE91ytoJpEctXETXNcFN0Cqmov08FbaLUVFz
cZEk5Q+B4O+Tv6nNaWuYLEOlGOQ/lty4ors4XtWQmVOIyy8YJiA6cWugSzRc1+TB
ZP1yiVN70q6TqflwClzAHq2GVsq2Z+TfscsE7H+XnmmlisOzex8f0TGFmneBYCwy
805D/w1SFR7DrsKkC/uvA5Bo05OQnYp63Sw6W/sQsgbzLxluuZoo3z/d1SfeGZeU
v/dl1jGjLYcvY9xCTsS8UPZnnHqt6mLUNm2asvTdxHW0QjGhX2WwOhb4YHopijBw
MBIY8I769v7IQ3//pUzR4j5Se6gJWHa66k3AIwjXhkyZXe48rBlBHjUHawkzgH+C
DucOEYDmVe8EefMHSAeYRIIlahL+U/2FTMhJfakgPNPObsx72wt34UwHuBm4L1D+
GbUeC0pyUldXE8x5UVq6RxO9K/AZMJf38ywIxd2f9W1Px1oGbJm+clXxGHt46YoF
zB1Ek2sB9PFoEnKHiKJ6E4yTRdTXVuyHvb+itLr8IJ9mvXg89jiAZuZLc97LFwJy
x/MWzNig2AmRWlvtPB0oU+uCLYoD9w1roKiDJCpVI/Yw0DwSMMgl69yGXWgd1Kio
n2lwITaa9b1k50jPOEXjmoOJ7uKfjUpM9VfQ2b/Q3OjsD1mS1DGj4mTLow5cJiwy
URuJuTx9tezVcVxlCCrrGmyT0n9E3FJRi7zNckiPiC6fP6mDRsicbXC+d52RvVwv
4SnATSR7/tvESK//1Uual3MiDvm216hGenWSZI3M5NiMyvfcMeYpgM/gbv+2JP5V
EKK/qZMVPNJIBM+YEgQP6DgpCx03Q/YVdeIzoYzJ7ZHMqOe56aokdGIShyZ1m4EB
Df5gSYEYBLnodvi/UZj6Oui8n2qVUGma95/NwHCUgT0ClwLdPs3WDMKl6gboZIz0
lG3rSsnmj4okw5zB5ZcvbmQzSvIe73yhdeIjwdy8KieF/+rcAqH5g2T7Vk5zBLpb
JoP+hrjcgasMyfoOyMc+0suqG4qu0WitLn/wAJvFO3WL8Z2LDNKddIecwDZYD16s
i7y3kdLGjibTUIV0fOPjqbkK7Pl/eMHuRN+nYl8WEei20q+hYOutEFsaE0A7EwPT
d29graZ4tB+3fg7RW4UkNpTXJi/Bj/leCa+mXaEyYOOlVxL9nYBXqfKkSCYk1sEn
lFpiTAh/cJBeXXWIR2XEWQc7NQb1qgVjZMCSK/gjx6ui458OM9o5hfjrQVimO8YW
+DXC3BYOp7aqQ67Let+wRoYjNd5pH5xpGOWRc/NHAYBvTX1JWFdGDfEgUv8gPAX2
oYmzF07JkHVhyIBYjPJIaT105MqJza7MceRTLpFvvDSewk2QmUe1V43yuWMaBOuc
k/dDNfz5t7db7ya1LidGEEYAVNFuPFKC1zZc3z8t+1Ccakle6UmZ3NMIm00Z2xsr
AJMOQTue9w5meec72s5VXsDo0+2CXvqLIoZvZ6uRa56T++2uoq78/gGBRo16UzAB
WJB9iZEFI25/BqrjE5Qg1gR0l9wyPCXrDmFr3VB0Zva/aw5yXjlM6rPyUZdhUm/2
/1FnL/DULI8uFpStX75o81f3Thdefq4g7kXzkqpvbRKDc+6S9xwYKImcMG+swoGW
cwRnzMsYuBAUlir9cpMlBRSDklZWzTeOMAd/GEsdmZe6masSxT6HEQgxdyBCfrt4
HDm8Wno8ZEkwGGtqWyKyQAVzE8i9ZukzVhvoBYMUYM7iD3cBatV3to4AzNClxHLo
osubbMNJrTqe3P5h0tLbv9WhtSw+LiLh6YmyQnmPAYsDl+8rojcxLbrBoAOvduK9
2qmTiXMjDv92+HcGSk+JholGvfPtmb0hzNFPiXFykXtGQbs457QOP6XQUeQNtBMa
NNE7ExhIHDe76Y32sLzNTFv3SkTTlKpRXTL91WjgRpoZ38dosHk4Exp4RUvesCIW
nsR0FmVHiuaa+sSO2LcCOMNeSiaAMu4FemC5xSbwRnEnnzYibjUc0qE+Q+G+4tBB
t4Ao7igVb97/czgKM44fy2ox7r7lgU8l1868wTCZvjuP3TZhySjAM8+WBsNMe4+p
KhunFuylgNgTiYH48ve1USQWSQD9lNwLPCjxkIiDwhDx9dwG7662/9OQ/xc/aL+w
vpjqpdZ6pc3577V7ZzuBSPlu6jzE1Cbv95dBPEkVWTcozMFl1XstM5Eeas0Ws6Sd
VIUFPOQvOJb0nOH3jeYT32yQwjdpPLTMo0dpn/C0Kj3i/hM3DI6p8aVa8sg4Ftjh
d4EPW1ZN8olv6XH4u25mLfcKy3AUj9qrCsDCJZzi7y1pya4vrXibxcQDVTmneZrE
kh585K7OmmNCNS0PW1bCbm2kPJ8Ae0Qx5IeZbl9pOHo90SbidnOz26iUjlJqxEyW
l4weh6M8irAesZtWpOQcfuL/LLtiWFJQpGWpo4x0L89nO1Xtc9COM5sfyH75M8Cx
DqMYJ01/Oo9jwY6jMRttnkQeDkfagIxgavnARqqWBXnfWHyGGguL2HCmlxmqWgGi
NFfKpA5BAOfqKooLxTPVauVTzAiZebNh0TxFYUXZhbGNBX5N8q/S586rbm9b0UWk
EgZujBdgvAW+EoiOID2rTlnEzOMCrgNRko8TLcWkwG2ipyuWKAPeLG+c0gYYSvjv
YWd7ht0xtywhCWqEknMkoxaCLRYnvr4KPtHdiYQJP7S+PN5GRGq6Mf17A1pbL3xX
apJ+qt5EHPUAOQMFqZZjNn11PEqvROiRR3gX/y4dXK76OfjfX2Z0H5o9y2PwH+Sf
zQlEDL0anO5FsOz0g1/VORmKsvrkZWkgNkOaC9LzcvZGl8FpUb8kXhciH49rK8Yt
q2h26oTrgRx1Nthr5Z8wUE0IF1do+ab1cGUDN25UIuxwCXfmb4KwF8yWA74WGHg3
gcHWXoJpiisgEXdCgFkz3ODAIeoD9EplNbO4CrNPKdzH0AHM8QVTTlcU2SD70f1O
AQ1IlR3HYQKZr4jZ/9P9OwZG/cBSxzFyzRYucNkHD0+29beQDKVG9s2R7d2iapkg
UkMyWdUUtHBxzfR1PoefjEWc76hzkRhllipVUHJKubsUNXSmqTB9tBcDE3fSsGHy
ikZaRCH/xbv+lctgS6OT7JxNT5aKwTQc68g366Hw1hJSN2QVQjVjBxXHMnaLzNPr
USo62xFqNtDxLA7I1OspcLFSludaUpjxSfAcL10Dc5qaU8eG6a3hWRnsl+zlmvqS
5Srxx8pNlLReGQW79CMrjgRUpMgCd+FvgmDaV1M9Gmbl5mDCBahFoSyLApssfUs2
0LUlnuK+1tyDj96s+GsA/2Au/OAmxlJ50PwpOcBDL71UxkLaUaLyBr/Plr6L37GO
7LT3/n+8OKcoj/2G+jCa4ijaLOhV4FvXVZN1geJz/xLclfFPX2YOPDrWACgrKyR2
nUJfJhjZFsvRzbjbVrEQ2/xPiV2vvC7CIW9iUMUG1RXHCpJ0My0IePUuXPNNTlKw
ATGliT+r0dDZXHnP1kIwlcXraEqlEjVbJBNbwZ77q+nBtq3P9981Ufuzl6JP3h29
uWfMX7JoV03k5duwDE/IT/PBKn4e8mVDNErG3hKQdNKxpe6NngiJiVRDKh3AxWsR
PjNRf2ibJpFbrgg4/JdV5rWVPFdqrSaOWGWuM6WVPXR67zYTLlNX2NGBsFuUtj77
pCN0WVeQpuYTP5z7y/y3QKcFhkZe9Sn4KoHXbpvt7hHSwilfFuPT9awdwXVHG7/o
3yW/i2LLXWw1KUsunh+Qy6nWNHmoypKSe0k4AqCBhV/auhv/oRruBfxNiF4SvgTO
aPAqJ7aLQhRtXXwoOUZURkCyPFw9rhpmuXuKlSYi4md2nUt08Zb0Geftm8fGjhUL
FUgxzDr2UESTeZwxhSOeUv7q/AAw+uvhb1NR3rWeFta2FTHHZKTB8uZukqpLJrWl
CQc3q/1hCiKYMbLsirLfawhptgwRwtgEbZS3yzcDQ75eV22gvTyJ0XstixM+pWdC
cH709drSPg1in8n86Bji0QX7Hl5LmVgbSamW1GN2W7LSNOA+bi4sM03QkanN5FML
bx2OhegL1lCDk4+0zm3tnHTsEbschHvwjcW4vmi6RyltkD5Hmz4iowdJ7MJaE2C0
dHRpYwXpptMRrd7Sz6UoCgZOOPwx3ke8Js7RgiRTt0PsKmjPK5MxcxMARBloklpq
N1YrhqLDbyqPUmRgkQhzJ+SQOAS10crbK8biciaCMY80ywheHUSNsdGIpi+bj/oO
/971vJZ+h3Jr6ZYF/U/t+XF57xpnOg0AbeecFFokQvbLaNeTfz54KUbLYRF0D6sg
HJpQ5LWOzxYZ2wvLHhqWU6TDJgJQ0ujNgKO8g7W94paXaIc6nwwujVMw1kJUac+H
EpPQdZH9McUSlgkQzWC7L3olSTL0Cjc2GZTmd+Z1YhUdJnaK+fTVwQmcWrwDMu0G
8ski+ZN0rBLUulCPAl4Sy5XWGik1qaVTX2SRauMhrlL/Y/HNd3GfJCF3jTiQthQG
DlsCzMKsspjGVQRTKTu3mKpHwekwLMaF8nzCRfszYO2Mc4MAQ2DS8lD7yRKYBYMY
6JRab4NqeUfyppp01Y9tSdFoSNJSM4wPJyL8B+WJYzILtAxX1uVBM21ZHg1RsCSu
BGBMOACx3qkwi52WM8jXrEBYN1acIP8qU06co4OMhC97+9V+kqL6E4ElpwvRe+An
mE7918k3niZQSz4PL3pqAhdPmL0E5xu4p1VP8tlKWEyoFUGIUBKA2ekS/648UA9Z
3bpXJBQjEFO21PhQQ8zVao6mnjxJ5jMhQrQz/z1J7SGpSsjRaMoipadzUbPsPedP
oJ82zVxHfFiuS41uHr6ZudkPulZLa8o1MU9s1fGq9trRiMJ+2ekUtwrtL510jlxB
EcmrxXUv3apnmVa/FwG8zJ6vQp8ZFoil5+YeVO/ROxstuFPT4E718aL0fwF2jSkm
l1RgXU8POJzh7yHyPFIvDPlOPmD5rZ9e1uNT1TfkumSJhktQx1AcZmmOjUd+K7d8
v4zQMqrlByU7PPlv9FakOd0TNUlKNrh3EXnWm68d+23Ks2uwp02PQWebodZ17lWU
/l0vqHEnjONgLcWXYLvL2J/W9ozpDq6EfK7JLRSmBM/sIKiycA9ko/mV0ceyGe8s
bSUTa/eBj++tKj44udVj5ayQ5tICpAKL5gQpf43dJt0p34GQIACFMsjfDDoa1YZ5
zK+MdYHr3vPZuoIqhlJ0/gzNO/Y0qlN+4EyDwfljGXI3UuR/wFKliEaB4pDT1v8J
n/yEkzBAhmzpqIPoMNrmLyHReUCIm2wVJcGDseh0z2IhQ9OiroSUzzLpiPSPpcPi
mtfDeh0VDxoiKUnOpSNQgTYkUr6uIM4kvIR3ZEs5JmY5kU8kT66baa5ZXkKbpvkn
M5QmTsYZHG52tsUqJhAcbyGJ0LF/DJFxwNB2Pb8p2G/WzeYPv6mHkpWsGNBSmDyG
poYLMz9FNz0Fw2ei5i/4IWwnDJz2RaIrhgRzj632pVKz3FFxsfTVdJF0/cip1UTo
o8oQntzfLor04lS1GwNX7AhZZlJcKJsRc/2ivAtK5kerDjGUwhbW5qg0dprqRO9C
KxwZTAdde9/zf6dAorgQXmw3RpLw6CX/5Pik2xR3Le41rHg2q3nOsBGgxqkhQ2fd
O8JBvAEVVJ1Js2ldGLZ5cy6KGrjQjQz99b80Dn02Z9U3Hut9z33YBRs3uLk/ZYAd
hnCgx/0fV8eXRipuQMV5HdIz1zcsitGVNYuAjsC2QNE0AhLsUJmxoPSfJ76GumSL
cUt1JLN9EJZNXxJKm8vZkAeO/IxqCRhuaNTAWDjUPv6h109KUaurHWBbDqElIhIq
1EN9bsiUw/ns2vyTExH/gR2E0s9XHwEIBh5PHEqQuO1KPnvR+vdziZNiaszJvRjd
DC+LXElU+7hfKs2i32OYicKpHXqg1YNhrZXN9adCRNfSPWSltOs5Bj+CXhfXLEzD
wIEHR9fVKL/8vP8TeiP5LH6w+KuuuEmLNCjvkTNHkVoZXxTbpW01BGU9h7BZ0zxb
+uYDFyeWGF87ZoTJLBkP3ddfmsoaO/2kveFGcldbGMfpexRuud9WBA0eog48L6h1
1Jx4GoBRIOaI6m7vVZPID5urSQhgmes+z8dGY3bK4fcYle6ozEWcizvG2E4w7uiW
n6g6hXBo3ML4PqNXoAcPWs45WIlsexvvI5RrMVWVEgi1dlBCkRpf99ET8j+YxrEP
6c45GcG4j2elTCp+3RPYV9RELXnTENoUnSdxRMQ6GrFRsD/IvFj2M1H7kXcXC56t
Tyyhy4VdvqfQApQXY/NC1x7A0q/51ATC48uuQSSlNZiHmTqYy/B9tcvKYWQEVhXl
XGoDEtcHr+R61wsDW1NeH+ycpkwXhkYj8/RuDdyzHmvgNqZPX8Wdy1VN0UxYrx/C
f2Y79Hylv3awBwI16mkng0lWDZlcyKDQfFGLSztM9s8iZ1NdpU38anMG8+wa7Dm3
+vCQYt4M7rxGIVz2WMSEUdd1VujzIGJUFOAgMqmBauLbJBzjhPugX736kbzSBlk0
IXrkVMNdVaApXgLXoN4YQPV5IIUs/Uac45ue0EicSz4ODRsAYhPy6nmlETGKRQoV
0mZcySEzJg54uIFTpcPN1w4e+HhbeSEhfAOdV1rjICYtXnFaXRSOatX394dSowlg
SqeF1Q95aRw/l26wKApzOLv0aRf+Hr8IU6iOiAlNAhSdDNL1/4Gc4D+6N5HO0LuZ
fSh/LqrslyIvacpB3TJL2w5fFqv+IPcZdwmRtLup85ywNWJejj/8QdmgTscoePtL
RptB09d90k2Lo6dPAUb+6Rf4eBcGUa/26OAR/qen5BO6jxTDElUQ69Uurs3+vzcN
NW2ltqQ7b17McxK8AtHf3rLEvRImwQsFyGSzh+I/z88QmZOUJq5OHiZW6BK8qNoz
QckULaJ62S5DokLa9e/YomERBRhQLT/tD+e3zaUw9wBQHuwKMDqHaZrexDu+7qM4
wl55fYYthRSEwh5qmQZagOJnvuyMj3waqdUXZpODhwWIdEf3+iJoebWCPsG/jRJh
KlxvcuIVPGpmJ8EqaPQt5QPpietc92aCDVSTiU09nhmfOxvTO+Bqab35R0P3oH1T
8KMJmvR/SdTJ0BnAJK10peklBk2OV38ID1uL4+g0BMHa/ZBigyMkXmN7pReinDYB
4epHA1ieA+H0hZEI4AUgXXQ21jRgI3S4wIse7MDhUU64xfywpvn/FO0Mjka2hb7X
A+lg4D5lRsYF6uPrKKVyUdgbqbnV9GYfdsJ5cucyJGfXaGyf+RY85U6kOUQ4ElF3
EXdbtUrP9aydU+R3BWWtnTHLfAWzkV4inVT+RmY165LcikUX4Dh1oLBju47207yb
4/CyZWGi8WwUEy7fKdyaLLxHbCT1EHza4j6rNRYS2EJQI1sztRr8ilgPyt/o3ZB7
9U6o/h67wZTRZw7svtCVtUAV0VIkD4fPXD7OOR12I39K9ewbZo/GbpZlKyMMPeL4
vDklJBXGFJ1ZBNPgcrZ9qJTjDrhCR3K0XgEyDMSUGouBxEAz61zt6qFuNH3I3I3H
8cdxn3gHOIMQY8CuGjKdOmgQG+V+zd7fyhO6p3LL4pLiH58N21b/IlHKR/fmV0+3
HPDRVJPapj9VdNyq5lZUhj1Go6Fmr6zgozsThKubWuEBms0WeBbcotjyGf3HKBrp
UbjFezg1qqSF3rZtlAul+8e1qkiGdElLybv8oCyQbeAqRyt13R424Xct2fNWKtla
DG9b/HAE4mkXYvexOWjkxz3O9LSX1PN01QOuCPhwUthqWNZsLPzxNwiwFSY1k8AF
FRfGvHQP3kooqD06pxdMnmJsr3u2TfLOThCIoSBhGfIzyrF98ZQP9rBEDeAbiYSC
LtpOXA+NmWqNneV10mFxOPAGIc9mB/mujYmEw5we6GbEc5GoS7wfAZAVlUN2WMj8
1VAqFjeqX8NFV/4Crg21xd8yzkbXdoBvQysI0sWVtrcr3K2rpYc3cwwB7RXVeOrM
/gUYkSiVvNeBqwdDgt1ID15AcOLgZNJ0tCrOBBHzzamuVzBNWND92o8CeyICL1SA
5ISYSi1eAyOPb18DkFLfpKtEP/+c0+YpUUP6PD5F/Nzsnsuaz5vcVef9cdSD60qS
jayC44HOKihwgs1EvkEa50y1jmiR9IpOSTlKnlcKc0Zw20gS9OwuFgGVRHXiWTlm
uVCMGT7qEaya1gSgXsfep0EocO9YV377zTPiCg3O+5LbbN1PZD2stm84k2+CF/IK
J9PGf0v5BGkRkgOw0wIUHrOHP7JlU3+MCXCBxkpt6rr9HbgsfDamo/GgOHYVG6nJ
yeMglbp/oZLtpFoDYNOoXuh18ubN/dqBJaAsQvSx2aK1ws6cr3aQKvi6LBYH0qr8
v/nEkxanOvNSYDEWT4uHm5IHbDuHzMlnqz+6qrVNeC50Bzxx4ksafrSAVvI3cJoU
xwbKytMk6zbeaRM/uXtNxXfWD/G/zcBRcqu5bHYOqsC7RniWJMSiVBsDFemcODZh
6C/q/2nt7mfOJNxveWh7vrGktj1C55UObTcA1rsDlFXkUlseXKuSZBsl/78M35m7
s4epCOsXQ5Vkq3W5h55udlO7Pq2459Hagz6fXn5NseNHOSn9Xf3FwCQZ159kAtiM
aByg5HU4tU/CJUnI4tP0a06yO1bgzKOw48XUQzQC8SpBaf00OFJJ8Ox1/+Xwn/ni
MVDDcYTbI47Oqum68+WVLAmFP37SlkRvJpizFUlDY+70Xeq02/p1e1HS9mKVsgmO
DX/HtOmDoM4VnI+AKEsfw3Ewk1U9z5POEI+ceuloWIIui8YqinVAtD5VISYKLF3+
yjA6D3mOfCCMNoV8yirGerTYQLnJSLJLWQWKLwhos9BWpfcM0Oc+4+HLZObiQiHm
xEoOuWo0NpcHdEU51mdE2lJsQ3NDSkMzLlpzGEcirTIbx8kDV3ND3wYa8YCtbF9U
0f2cAL6HAb7OtxqJUjKxV0fWa0w+n3lQdfMOAf4Y5JcKxExHRY4raivPw6qIFrrr
k8hCmhHmy/7emSZuPTPnem96LXPFW0ojofDMPRYqOA3rXOMhbLbk2q5deU7i66ss
N962ehjWI/TKAZ0TPgZ8X2RlKORtVhkXc3s4tmrHAdTjkZPXCXQvKIyVCGfFF3Ll
7eDLMBvr/KghCZCRcVxKw5OcqlN8jkq9yG3kw+vpXLIteEEbppxiXqWc4vQlhujJ
bPBlDJO2oac759EoW2KPni3oZjmX0Yc0gZ7CeMGgCFncyDBpzqPKZF39J8iECTya
3RkqSnxf50AyUN7z65jfFCHDbL8YotgSHFMYBKerqWMC6s6VkP0jkc/klJAbaNWD
hSDP1tLyAQHWw6Yqgv7G5HOyNry0mNHkjAoFkdTnkwZArL1pNt5fidkmUJbNA7fB
oP7X9c9j7PruxEH/RzH26HHxhakBzHRjjZryDcKr1dgLXMaBpIqdjVoedmDeBCBg
ZYHCkFrDACyHo7lELFdnQP78exQSCZiSDBEfiFSErQ9aPgZ9e89GIAGbi0LC3PKi
y+0/B6Z4SKpUgEEzaiNDElB8Ohm565Z0YEjj5EYgNsn1D8iGmm/ZNqPAD2HTIIFJ
RBpoX754ZF8UOEt2MmI0vcGa4zOVo47zRQaFqRnXlOnr3Wctx+m/5rLYVIYk4M5n
9/erWQ71D2JZOX12bpBhORipD54V3DBGILhRf7PaqFbG8tDFzb0SHEO89iZ+byJZ
+B0dEYf5+MQNqWKW+KXXtqguBmTYXhsidgcYMPG129Jo3pAEcasG3QjwDUKjC6M5
CvvzweqAN5ytqZa4ch+jPmLvEHgxaETpvgU3DT4y5UeNLeiiN9RwppXNhB/71Mov
FRXOKWDOBBY7i/ihVMzP9jSoALlMezhqwimsvcnQOf+L6uG6esSvKg+bznICZOdo
FNZntmoHZJ3x53YTB/5ESLPLTFkUKLjUQ1xI3uzL2cZbXwa/7CIULnJa6BLz05nh
uL4/1FERY6A4SPg0C8P/CoPdAyBEExTAqIbPjKBq8xUwqNZygDCUb+85TSX44dd8
3BKrlbiy2jVFBXO2jmdf31Xg4AME0qQsz3FeAKSXcTzchZqg0R27Is+aYav65xGg
3hzCNKaF3tj4qY8OxIjkoT8lhm1BtZYfDgXD1OijYV7lYFp3WzvU2ZDGoAgRLzue
ql/oOjMA2OEb5S/WZ4EOenJ4VXdHeSbfPAKFh9YzN2Mvw2nR2JfYWbuK87odUwH5
QCDxSxkGgEKJfBjys7vvCH32NaGFawpPkUK4eYmcmSMdOdGWGl58VaDDQgADGiYs
9gFh3MANHWW1BtSZTDa/KJGR9M8luTu5BbZ9ecDUf8Boip9NBI4I9SsKiyevtNyc
Yrx/3YsyTYMC7gDAJUwof7eI+ZodTCUPOlac9eqaW+bUH4EDLOp/Tr9QT7oXaM4O
jTVU6SP1kvymGvIvoSMTuoWC1aVl8CnCS8KJQ3P8ll8K7GC1aGAXCRCz/Nd2TnaY
YACjaUAlfmDCljEJ4pQ5iDHOOVY4qQAjmY4gln1SV0WUO8De4TnU98ohNlnzvo70
YD0i4AV2UQhcGztHCetC/0Vs9+2NrpHfDi1eytdRmk4Tq5+eGv625ETLehcds80C
6+16YqW9wukT/s/LFI67ge6+oCW//6wwaql+SxeW6XQkrGtVK4niqBhEtR0YzlH6
lRTTjW+O6uoePPs38JH6kLNMXnaDSNpmZe3W61D9EHgDhjlYIXvLxQOAX/h0LI3F
hjW716/J+ohPGcEZQK8jNy/8p+SFWIdzRrQeQ2J41kmc/mIQHNaASrGNVi71NO9y
x1wrEEBqDTVU8CASDUfanhzHyPN9hB13W1yojagFWXbykYEKfbLaOsz0Lt/7T2/q
wQzHsp6FUXsKwUiIh1dxP8WEiZkRkudCux6E/g/XUFy4eW4wroWY7wZ4KE6kaaKl
C62EOF5GoegzjTJZIVyGw1Hg3n44fMxiVvw3goHBL6AQ8Mxo2I4EkM6x8mxXmvJH
gzQ5XrsicmK/ODFng3doPnnnnnnjgTaDUqD/Etjcbyt1JbITEctqq60+gt4ISzuH
7MNe4SubCcCQsxwEtzRkBNepmrlWVEOi7KALw/qPM1PQjOrbIAYMxBkJEnR8YEGr
UnM0lDye/M4Vo2v1sO0bHF+mbR6Bl3IFODBFET9aIcTH9kaLmnct3bTNLAZdpYT1
NOWypdkD+IU5ltDYq6lorKFchcS17wvbC8ZaM0ltZXDhMmjGnrEqYfnODYW/MkBg
Zxqr4n7F+0stY8zgGWXdGswOW8BrRlDmkITa54rOkwnbg90dWll32Tmk3txPial2
Zv2QoOFo5pklCizzZS3oeuP3wYslFlryrbyXyEBAzglacFaOwevqqZ6KmAKeCNZb
Ey6pgqn6Xy0akxyt5l9SEsd1Sao/IUWUC6mepK5J20s4jJA4M6/Y99XPgLsVxlQf
vMpgDrQDooQuWq/7hhDDMc/+yt8X9t+3Bgzo65ymdOjrJIm7UkHMgLhNItS+c2XB
Di2jlyTuO6pBePGrtFk5uwrg8aVE0xzWckPnwmYn8UM/ChVAClUukfTC/STOleYI
eQO27cvg7eVGnu194xXRrZTdgpigdm6ir/hQcsSpRDGawx+qkdCzdlrsLaTOhvWV
FKoQFKw782Y/8+nprIMg1CcBh24u45RCMfUAAqtDuCzSvPA5o2z4bh3mOxWwl4jG
UqXfsG3jfy6fslx+oH5kO4vye1u06VsZUjBWYqswHP7hMIcichER0SDv5SxXskgP
JfXyYPmAGoM0Yg9yAZBzDYVYd0A5DWKlvUtQp6PWvmribqbbMAJXnK4EtjKlwjb0
uWSTgK/1sj8PcQaxV/HHgKEadpLEtjDbal9bIIPweXY2AqTLtk9XNpewZK4w8+Y5
4VA06sXZkghHeUz1k8JN8z9mE2raktgGq6Zpmdn8L/R6rwHmdptq9hWh/LdmHnZk
tQyXfJ3Uc0y4AVwC2+6OBGRr98Pu4Glla9zTSKQCO2/rBAmypj3vDoapRlTpIDjh
rSpE3wHTPgv+cJNfvBvFL2biAeR1dZ1r1blL3D2W2eOpnt7wIJ0NElK1oAKZ+dJR
e7RTFl6W3LhbzwKSGYdADqEIc26tgRU0r+VcjTEdvsmXCSBi4aImM+5ZyeT5bVc4
watJ2XU+5ryxMAHmc47tFm0r2FGU91pNCRbGQb7uu7Bd3F4uz49c8F1FmuYBZiFJ
AH2gI0U6cjWQQ+3k1pL+A50QWeF4E0hh4EZpDZsB5740IuAn5s91r2Ri5sKlWX2/
IjqpD1YXVhiVGFoh+SCbe/r/nN7+Csqq/NXJKjhnJXyRbHaTZh31j0hJSqzJ07ri
KCr9qubWo7R3zsZ9F3qGXQgXrd+0ojwiDIKFAmf+3ZGYUjEsn/6U1DboZ4LPFi6b
SExXSEJoKDLYSF6YaaddoezRfFSRObxHiUEIncBKRed7b5m06o/xDSrCgJk35JeJ
00xN0ktoplPRnN2osjEL1BkHkoMAQT+zvJZ9aim2OlW5JyRWUndjvm0qsiJwxhGp
5A/XIX8l2jo69Pz9+icEn+Ikh3QA+9k3DCvwBRMt1MqM1hxy9YyAJngCCK+l4W/M
Y7QlBBTYj+Mu89yI88pO++hRQlQZ+ekhgQP5C2dfGN4ww0qXgp2SehFpg1QY7RN1
ZXrI9xobydqLJvWladqbvj/xLayZQTHwTQ/H7qEcJ01j4Ibe9pNCtivKQUFO6ah8
cP2RNkv4lYOfq3XSEJzR6/QUI84dUHUo5t693HyW7kAfKIeXYHMwUu0I3Hf+BuNq
Kg6LROlpSW9NJL8iUO/HpWoCZJhrQfpPieK0vvRA+GVFCyleu1P5poQhKRs0Yfx1
ZTBL7kDPaceEkaubKVLawoXQq6uS2LCt7NSXMBNXFJEk5DrDuL69HvPx/hE3IL5j
GIFKOMr7W/7hiOsZ5JhKB0yNqrh9Wy+7H8Km4x9/mjZERGD5B5itOe3/C/wZo2IB
mG2gIYwXTpcX19RvFh2tqMO36+gsfxaVEsJJFVqKB/sPfvevgihyJU6YZorbHD3V
UnB7NUiF4sP2tDhWKeXYglP44fT9CSgFOpcakEy6GAeBVKydu1vTv2xhMKWJ1oJ2
Gos1EdOSK0PdExaxGW64LK5jEyP1yQkZBltlig2ptZKtXvmpa3hI1cFz/up4NqV5
xbA7NeDWtDxAz0nBiwGZXT7vz8WhnV8tdYJhSq3kl5JniBG3T5sxJaqtEdzqkmKO
fpWIe94D/wnuqQjjXeFJ+zAc2TxUDe9RpwcqjlGkVJwwwXwSCF6bW5+ZqqqjGNyW
IZf2ONnO5ygbiyr5NLpQs1k52pHkEUVwxPjPIA4Ay/8H2XPYzrdD/U53qD8/3pH2
NgS2FMc6gEyOU5FyZJQqxHcGPo3oQ3b3GtTyxn1sStiHL8EIETlR/TAyDontdIsA
n3JtziLb1CEQQEzXBO163YJMXDr/T0FMH5C2RcAO7CRynbplTzq1p8HN0oAEytwS
cPJy+qpZNeYftG5iGIj/Q+Tb6QDuSY55hI62XJ6zvVaV463I5qhG/OUsgsTqqefp
LPHO+imdKUvkQEXoPMauXxhO60zsApGrA16XFRALGLHIh5Bl5a0C4DD1T2AxJj6B
nNDWWC4VPwju5wlyBk6XZyXl4MxYpSI78LTQq0SgcTmuyWYqGF+/Cinfnbn8XdNC
Qkkg567BJKPnTIVX85IGlNmIjX/iJDXgQtil5+KNQ/zILf5jAcdejh89lunEkVNj
50VTeJxWuuEeEd+nXBjecrnkRgHPgf9Rk/jyAnVe3CguZp2PSvCwsM4lrZafxIdj
efboQmqcDpjXtuTSsZpp9lw+jHOIC0uVYMclIuXHs3Yfd9wOLbbNbp50oOMy95Md
UqTnNsEqwoD9uJ+wV7Cc5Vfz+7mVOYSV+2vLhtblJR7CAy7qpS80bSyRiLoTfUqY
vnhpiDQaGJf2NUXTmY7vAP08v3xsawYlatFTgcLpIal1aZrQaCAYCFf8eDQfKlsh
g8V4JTWMSCKadnfPbPTkZL5TEbeqZ94IKPhZ1WX14F0cg/pYlOJK3S4j6xh4gPmW
l74Je3DwDSxIiz5Fx9C4JxZ6/h9DUuqt5YcmLXy9elnlg7mwFTwy1ObQmE/YIwtx
M2Wt1MpP3Zs8amqEm56J0azkd5zo8eT2Bkrp+nSkEKFOmAXcYvRx6MdeVdGrGaF6
oEefcwNItbSJXkpHneB5S+0ipL95pL0eUJbaNiFL5eR2/Cq/AWn0gSsDKBQ9fjp1
nyJxhf97dc2FyVQqzUKgzKXq2jxNo6782dDKbxelEoVnMJ7ZzXjpEG5u24zOn1A4
pnOu4IW/uCreTSEzOTc2Xe3gDqT1sHvB/OrNS9KcKezN3bvPzFAVC6HIBUDzqXu8
VCpeKyhlMNtV3Ng6Xb96EbU0xUnPchO51oZPnnZ9AB7SIqMwlDGOu1uMKIdkOTLZ
/PQPh9uXaNs5dzbZskEXXAYc7UhhTbj1470B3TWWeAFJYyi/4pejZABbmYz28WQE
MRWf73UsUZcGgyzirNzZySbfwvSN8p3vqj6U6tM8TtDvwmFOpRPCThrGkGGVUPfL
IUnH2TDbfk3eI3TIpbKp4RcVTIQdFncul2gGqy4uM9y2l+CvgYxzei3kFtCZtgFA
Tu802K9C77glRdPsZgb6YcA5pnFvNW+swghkD6EKelRJb52iBBrk79zKEHcXpbVd
Kdpk3cB+aVmC7MGGyQGKmgGBX/QfMiVWCe2sGAmR3sSkNex46uk79Pjlk9pS4lBQ
s2jYoRYdGrYZne5KY2ZDJ+B6rgnqMh+KuCCJJ5t1AMfIQ37lHiIXOJJ+lZAD4mI3
9Z8JoqWC8V+yqXMoyM0Wlof30IXbgRthboXENCcXU2fxbEzYFd7DPTuz/UmaAJOb
msYnzFMC8vRRNFYrI3Cp9lppLVxsBetyAo8ThrcZOQ3PtwKN2ItyVUUyEPo5T5pS
3gAxuylJ/25UzYlQTD3LV4Ea7ZWKkvkevdaDUHdXoLIc0pfYG1Jbpe+a0QK0in1q
YgPz6ccbxSatO54GupAUCcJty783wuFeHj0DssdNVdms/806PdPgQIE7WTS0G33G
95XHry/xLlJ1f621cp7j2RAn3JYUcj2VJ022MGQmKoVAln6GIbwbI7e6WRMroNjd
0ASizkxLm2P4wHakpMYDOJVaIUmJi8W3d/4Noh00ZHj864iaP2gOzNGdqbRoQN+z
vdmnvGIEziRsb/KnbfvKmC3t30yFSq86UVRiLsOFWiKl3cc4dYTyQxtXmu0hc6KO
jIU6ym7pKhJh7p8KCHLR0FoEGS+Gp0jO8es5KavZtoQmME1nRV8XdqS/UeqbIzZQ
GoiNAVdbz7UaSwYSmuEoU0P01AT7Ar1T6mXNRZdfH2IHhyRgc3rMsOfydYMmkFCf
HG16zB1AHUQld696EMO5sJ+a1bUzu0uCuFRnzRV77J3jAkau46njloT2toTmjcAv
mwnseIfAAHmFouWFZJqMmBmvunrK7Zwt9YIuZfJWrs5xQhIEU0vR2XyqLf8antvi
sRDQGEmCCbKjfOJZ4S5DDVXrD99xQzUhJYXVKWIixaREFzX/bXy0auLCENq6zQzP
NBX6SzrTXr55G9Yxnp2fTG6zElXXx+qId4s6GIhYDHgG9IsJ4yJWkPoD1fnt2w0d
3R5tCRjGL4mC9LECDBrgGhkJCIvh7WWvnXi+0/z7Ra/7oF8Wow5c3BIGuItn4ifz
2++N8z/B1SqFDTL9Hlpd6MKk/m+etlD/2tyKmIPV5AEODPS1QaOIRHct92NhB36h
ndcaLWSf2+hP6Iihru3YsyU9gRP6qvzwjr/YHvBU4BWE1CZ/hsBUyilhVsypGqeG
BunXgE4ap5kKxbSTMVUWQCxQX/7ofhR6pVp6liHJbYrJFtQXb7LTUUYfqupTtqIC
PKIsDPv9qWGf9ytXYQ8xQiTDJfG/WGcBPblHIyE/UnZgulMyAdic0ikr7jWE7yJy
HR4kQC+mPGBU4YFXUWegOg8YbcUZ4PyAPU8psl8qWjfDvOf+wKKLR2KU8IrlfVXn
uFaySh/RhgtyQfGz3+WUnL40+cwS4fwyk0OGQShtFG1WhamhBcdXSZ6W49egj3Me
DP9dsm8kM8DyxZbPP3hdttJat6a6nSZcBZS5SL2Lnf/zWnZyIEubxFG51GoPXArq
IGqtDqAQSUzNjrlH465l4/7th5Ydpb18r4gJol0inRICwFDxbzL4IIlfd4VY0i02
9RQW75rIet9YUuCCVob2g3ehqqagprSDlj9bl2Wq6EYk2+wtmO7/1DwcjilHuz3v
UbZfkcQ0i4vAWDYxNIkYMcUVJfPjqGE3JXXlZFh+wnVHPPuRvqyUQ3pdbCXKF3gG
2Gxs9kt80Hccz6ZgDxNG5guyESYHhexAC9RRlxkL8oOvul8MjZYZ+KTRiItdSkqN
HhrAZWiheXFkpmNfwUHi4Z7hyh9vus3dsZWzMTkwawFPBzb40/IHqgeHPFlf1Whd
Z4p0IvY7ZqWOucb0g9gircFRzMhRSXTQE9XOWp2UHTuJF/lR9yuVuxrNyiHp2CE7
k3xvXdFPvN4eyx1kaFR0/i4qSgC/CXN0PP9TgLRAeVAM+hY7bbhMZqoea0xQudkC
uro51P1Iqn7eUA9FFO9viWVDONrzt72T+l3/18zuA5BrOEXyx7uIFASO+Oo2Zfnq
fFPuAK7kaiD4wzsblRbY7DWVGG/KQl36x5TxbupviBVowuHru5nopnh+aAuQvwPF
vPFnBAhYd9Y0Fa6c2lipB5P3dWc7KsTtOv2kdEdEoqg7mz3CxKyb9ubhX/6uP1PT
vUeaUuJzqRG7coecp6xAujB8RBPYcXSJOq+m7hZVQgBpYkuiGYhTRm8qAepNFaA2
EGTsmn0QI6rsqgoagd+9McWkfLt7tSXvD6oy4jncDNbnsjBKDH2RIkFtoPnwnuh5
ZMODBJLsK5yDuRtyrzspm+iUyaDabv7ik8RJEGUbAMEBSAGmnPlkh4geCxCdDPNV
ItA+RogHtT5ECZAtFDBP3mYnPujkYWIalRlBQXBnbW1Nm6ryKPskV3mve40DLLvy
Ti8xj7dAJfB2p0a+2Kxflfdun7X+2arD9D4b5UKnGrzvnk6e3evmHi73U9oqVW43
1er9WOxaGS6NfFkZY8/5Z0DwIyHe1a+QXZldIQFEotlNI9D6tnNUyCjDkmxMx96Y
NPG5LiFsRQqDCDsnOnGZU3ye9zbN+OAGwmFhPddMNk3f7h8Jln2VLJrHrgRZ1YHQ
zm2vbW8LtNDZWYQqSmyQJN8tw/WXL+BYvOZxr8LQRrmaeFRxcV19UcaEXu/Tb45f
nVJBO4UxZf6ivgJfQGIw6wpheOGbxoG7oH0OcCiexl7ZjXCL2WiVT5xD3K80Owl7
kAAkUN2axH6fdRBxh7Iih2V1o+btmriVO/Gd/wgCqQble11plQ5Dsb4VOwlKBvI8
0I0ECQJPMoYm9jN63/bCfsxEP/O75p5Tp73CqOZb0ojKYtCw3lJtcJ0wZhfkiGC0
l0M/dIk5YP3eJ//hqIQE6Y5DDS90MPBU+A0BkghDrxvRtCcKIMdCUT4YnxnmnkFk
KnKU/l4nuPyBtCIb+54jN7ZzMMKtYONiKOx4XM8IsaTjNGpFjo0Duh5Pa/6/4p3h
+iMCwicqXOJeH68hXufH24rRSP24J9L9WhUqzfhv4XnRflNDRjU+XA4ggEyvtTD/
DnvnNzViNmp8pByqM8GGPZBSmqnpR4eu708OYY1TScZkkdEBE9xPcSSGVzJ9yVr0
3Ue5ElwVQ9fG6y+NbUuv9qSa/pfGtT9sQKHSVYOo+VfeKoras91hn1hk/ZXp+0cr
DKfzOEkUcMPELp6plCUk1voEmBLiLViob7D9E3xMeiywi/lkdwnDG5FZfbhxANgT
vcjw/FtVUM+tzqWzR9mt638H3ju8CQikxrdv3MD/lRkig9Fs3BbiaP21k81jEuIn
HEZnttbRgXUfONFA3Nb7TILenEaHqC9Rc6ajKoENz1/wWbAcDuiyyVG2qw9v0h3a
Ryb2Td7idQ9WFyBaEX8rdB4r0oUDR2gwTbhabdsc3rfud9QmnpwhihS9X5q1SNNq
Z8wuC1uuEFRkMtMfSC8NO5BaaKDg+2ntQ7N6LY6Hkwz/g72ls7br/QDtvtXNb22Z
sNBP/RjG1eBJLzDQ8Vo7ycBwfDoLgLIrKiaFCYSr2iiar8AJO1yqPe/AV6xQ4UO4
9eqpk5NwJ2+MimwKKEjlN2++wouACV0Wa63ubrGpY+eqKQgtuloJa0PvWRv4eoyf
peyBjyEbeGAkNcsFr4JCUrlQGuWKbU5R3jOpgqsz915Amrx5o6XlL2W9H5Ow3/qU
etgmLKp4TTNTMDfhH7Rl9o856ah4twwgWntqQ2OnbaZcJs5RVrH2ltgzRzkVxH82
/HHUYZaP2jjHLY8DdWBLFbddRGQrgj/nM+CWEePGUpzqktQcX46IH1KkmHrmwefp
Je+NQhEYqFyuP9i619584tDfFZZMRT7k1N5EXApn2DuS+ihtDuAOg4FJcfsp5D9q
dRcytWAU4qCUztMWeC+mDWbOh5PCYmofTXjYBwxtl8aBBT8yuhU8WAOfD4JmACAC
blL0FxdlUiuw3gs75YU/Gt7+4WD7YXU57DJ8p2V9n5Z6vVqBk917Xpm+HdPwFHve
S9XgEu+Ph/vufVop97f3XdS+FSb2h4JdoMlycO3GG4/7tvx3hm4z0WywLWRc8zKW
OIooSy+TLCz9tMc3PyTP6bx0Upv9qiwT7GQCZo3kkNnLjylYXG8Jve+Nb2e0iKpQ
YBxcJOYO8s3Xap4zL37tQAgPhftCp0LxT9yHsPocAsjzSDt6pzLqfEx5VUMO7iKD
UtT5XXNhl8rN8hn2nlkq90MMZDmT1eynK6Nk7U0vKuP8npJpwq4SSRIkyJu6TuIH
SoaD/0ywpLhcl8tVmoHcKyqiVK9vatAhZ3ob0iagM6WR5TW+gJRdj8/ek3eIPtVc
W5OjIT9c56nYcH6vRhhg7wu1YcZUXuJuIRxDN30EJLYLEkr+/25Qn1M1/AZ3FF+L
aNVwaYd4m4ZqNNSdbcrImDhBuhHwFmGqAzWFFMXmhCcpd3/DnYdoqvCQh0utBYce
iiW8iQipu+lFiGaM7gY5tR3aijVQx9FTHtNLO2Wy1cNfgoSzpLVCNyEQ8nz19UkX
mWZrgSIv3D15pzDGbpyS4W1z6uVNILEXuSxyRZcqwVDW9R/ev4/YquV2nkpy5itY
3iUTDeRSRVISouJ8+cMlILQ6Zv7sl3aCqaIKpjaRSbvSWBx5GdqaQnBBidPVtz6B
hZiodylLCxFwytUi/+mlV9swVgzOdYE04edCQRnC7NTlaaZmsroXQCsjBuhdcIFE
UuwP+jSNnwz2hgcepJ9PqcXyZ9OR0Z5G2XdcWyF4YnV/SN4Rbx5sEBZ9KssVNgJ4
0fjbbymSNEAwcN6jS9b0srVBrRojy/8v4rxh/pXwM9ey9kJGKrgQ0PWZ9+M+slmo
eKQlVFBsKUyiBSc38SaOMCDSIZNSHS8Z1rw1naMXJ5SpMzhy3trqBuTxSCArga92
xOkdI6BAqwANZ6vFgbhtUUqivQ8HhMqkULt1C8mbIya0MaazSbbPHFq5VBsdPvaq
ceyxQ1kDF/R1+knJRO2/L5aGvYEX/iQFifBfNXv9F28nLC/Mz7ogAQZDGCxXC9wo
os4kU1NWZSt2uZ+wtei7LYmkSAktCmqMQMoUZ7G5rtGwyw5lDrhNWUAQCaTgN+UK
zg6+buy/9GuuVHwTFSNTuhhSUJuTe7hCg21otJtjLFBiG3LoBYXH8Tn4oqhosPIe
aG8hYdhAHgdcN/2dtcXRDHIDHzFQWm75TtrHALPmMKPrr5W4x6DuBd+RTwlcmfKR
Fshl5qszXhUvgsn3xnoKWeH0gy+93Srck5yQHeZlIQfboVrOaBKaSIZ8L1vmGrca
ec00M6u611mVZfoWhMZ/N5GdrsMLzFwM3nsZ9wlrYZsjmsA/zGZKCwnuzFFQFddw
1WeccRIy3+xqaH5evStSNvcjOdH/ZWzqKU7w1TliBw957g0qyDsQywWUq6QK7XSj
6jRNMp5QxUaFtNKF5eEE7f/Y+GazKyZejPebf0R7Ta3uur+AxMSpohEgjt7Dm+r3
+JodcMS8uPrjn+kkyQiux/H3ks9TTP+/3kT0rCOov6Yzz2zfKzuU1tJ09hHLi8bW
YyZ3h44em0yI2quzFI9rnq/dARPnWLXv/kZBOvfWyGGEWiNk8kGBMOBxj5oVD2dU
b/z04kSt0cprzT+Dzy+LjgWcNVSoqGrkXCksTCpeLjZx3qtu4qjn4MKZFU3M9VWO
mlX0qOpF5td5A841npGiRLfdbjBWRrWLH15t83QL3rfrYc8u/U6wYjp4Cr3lXkLF
HdqEpv457jktvd+wjaz/LqE5+5kiWhIm8dWC3rb1pmoNBPRsbq0WFNjzCV8NPylR
tANCIwDa6nPAstWHNxGKedgxl58km7ejbxhXgOT9GJBwarMILKoXIqU7+By+0fzE
S38ajPg3h3aUOfhlg2tcXYhgJHicTctyqKtGVpw0riTmOBssWQTsduG8Nc7wOHKv
fDVOazltpD1iv2X/49Sq7xmiMaZ+Vt2Zs9+69N8JX5gK6vNZJ1JFHx3nN4ujZUHE
N1XtGaJ2yPeLOUHExDSRSSw9CZhJue0Skt8SxDvS3e+IOtO6kh5R7ilrLjKuEmnB
5AzhwPAuU8gRCIIvcgZaL5+VNcM4XYwKnJ90tH7f3Tnn+91sdO3Q1odNT8n/GDOb
MZq3YVwUEe22mDQNhs17zPBt8f9Y483K8AhGaQwilW+ANMap/TCY6N9VdTDM2d1o
rEpBLbaXXniHVU7Bb9xgx4xQcFaFYuvpx1ZTz/RvgVw2N4994FF8Y9dEgpPKpXSf
Ib/lM5YTDj0kFa2GcqYRsNQ/l54YyMDVLsj6vF8VxphZFcAOCK9cJM8dOXCDuBpu
eb6xt7JTcGL2MEBMQLBdNaDcleMmFANiNctFrNBYVygzge/93Ju6o+hFXYlL0WPb
UBKXjYIuq4IELpf8iwydvEg7FUJ/LcAPeGkfup7rlmKj9Mz3AyAxPfWbWJGQKJwa
nagsM1VxmR6T31pb4uVEEmD/cWAcfwhpXaeTW/iVSr3ndjmK7ZjD9PvIzS1wi34E
mr88W9ne6LSGsvRrFy9pqxoGOMU0BtISy6cIC+9lH3MxlZsB9KMoqqot3ZMJPErS
uHG5r4/h6olb46AcgtCafzOmvEjawJ72tYoMcz2n8ovlG95bENGL9xR0OJyKG8U9
tC+aWAqoaApq+QLII5NQdHu/XI9i8K6oCzFi8gOGA9zeYxqhSzSio4Ce70zjY8Nv
WvMhM5Q1+HEJW7E6XZFowJM20/OJ9ZGNp+RP0n/zvRVEW8tbS55kTypZJtZG4QJQ
QmJIHPQ3qrX79Djy09zOX0Z2CsK5ydwOTe9RlXwCnksPMqplReCtWq8oe55B5+Ac
wryyylTKnRN2kcGGfEbyOcURSX3/aCfbhXPNJlQomYYSapBLsQJPM6fcG45cvUDT
HJi6uiMQhNAmTjlK9U7fBDMSr48uO3FOERnvRYTEpYwp4HO21n2afzzCZI0CRwrr
IIl274krypcJKv28dtjN5NyPwn17NwW1VzRHejiAVsaegX+FlgdGCNilofAR1Acd
YhxSIYlIwg+et6XmtWW5Qdc38CBK+MwR37rdgH/WwaAkcSgzuI10wnyQlSOkYPRj
Ws1UHcRReXpOzhRiazmZ7z5xbB9KAoHStG1p7E+o6eRmLoLfrCvlSF0IMGyCSdCf
Hnyk1HnKFW4Ly4mcb4Oy54BA5QRic/LAa8YRiCxz85IApSXk/SSiTxX8VpPPr7AB
j79ihto3UPpf8ynr30mSZZRktJ6UMH9WgQFOH5VOng4AI8PNYQoXUTJ4DaM+QW33
Awz3iak449Ze8RSLOxHm6SbFlsfFqYtlSiYpIMfri186S808WR6PjNos9m5Gbips
H0cE+mO/5JzwoMBcvfvli0SCXxv2VrPx6qZbjFUOswgxlT09tM7eBLrk2PhC5eLP
iZP9Y2k5dwvuPpi7Y/8JmELhBwusCQUHeg76J+POjSYEu7dU/4UOgCUWCjTOH23b
s28g+hDEKG7SxV6446TQgnuqqji0YewAiz26G6ECkNjcuEOqyinf3T2P2N76MMB3
w8EEk/Rp7GZGIEY0hNTopNh6KG9yXOBR7Cd1jEFrB76uWR5CWOe648UZJmljpyTg
e8x9yPWVpNjsOLQvZOO2A0XPTucHu6gK7EAFsw8OjQ3MlbHPyaqG54UdMQP0ySfI
MSANjWW4lA0xuJju8FMeut3nmGfqDBQEj1PzFlsyptjAVdLOKFc6iDlulah4pCxr
fALVr+nCtebuScGnm/0SGwB1yyIfD7+adtQsk1yev4hz/PZ/Zh/ytWcwabfijk3I
4Fvnc6xXy2njWUths2SzZ9vY+MOnf0vLTudz7iXsYaz6D+lroWbK0POyDio+5qZ5
RuIF4cgUoisOJ/uVMh/j5n7ri4wIuxGRvSMP9Z6CXJsA0fwTY4vPBmDWO1WPwnzW
5WNawEotgfGwuMw637rVKbgyrWfuvBvJq2EjVSbGT+huWE6OEf6ZNpVzPvb34Uvw
6fV3XxmrHcW5oq4g6sFJf8R/2JDiIsCDYobHf5w37TdqS7J7TZJduycEzzf6Efky
a9bYFYpUWQQAlsCPdjqUq2bWK8qdEorLq103sx4rEzkhxe5xtGGYAqJCUx6OD3ld
hcBSmBoo9HRgwtXeHf8AjwgWILsHyTLQ94a4H05tvt4c0Ndm9bVIf7jTLTLgFOta
ODhppY8DPKU5DqgKtRMPFGGndiLXOUhza7iwTeHl+rTvG56ssLc5IY/DsLT5uxBQ
Z9hMv+JSBzRWFtPMJQBNeK1dCOvBpgzh3NbnC0Ejn2eK6wHvvu/j4hlTuu8q7Xx6
AdR5MYtZYkYDjgK5rBFLD/nX/NJfQt8+lMermcsPgFTwQMXQWUJOg2j23EgSBxac
jhgASkD6DhusC+8AQ4EV7knlmNlOyr6RyZRz/11zPNmF5u28+nulk+jFttTZFGVb
m6h4BEO0aHI/XhKk8WZ2OwnD7KBS9t4hVrwchSSQ3m4dNFYdiR5+qO9MvH93Yo0q
WAcE1YFoBZbMXQ+03VYenkSLePAogn5CoBpvhBswjCZoVIw0UVAzm/cBM1Oywo7B
evlOjaR5gbzGLmIyvkE1mAkTjTIoF4cip41WW4oF59GpVtVmxCWnMKlPLapA3Vx4
F3/CkXbMlXQWlphOJ/EnM6y/co3JS+ptk7mg217cp6ZjCRK99Y6Ih8v1wK+fFNkG
QwPriCNtDbpDbmvIl7/WrLGg5njppVd+JYLsbtZgJ7LiyIn4uEuxcdzRFmAuWlgr
Il33OKhwy1gz+IjbJ9qJ0es9napotOE5tH3oDnodSP1b4ADBSlhgQLUokXrG1g/p
oBjzxw8i8QMKTMEjxu+mzG3URUF0ZFn1XDSCLC0QgQ1x/rx2fwRDnLMImsD3+99X
hJmUVu+1coxg0XhmEB51P2XwLlnLiiyubl7Q0wCU5kSYUO5CBk9V4jsF5PA4eOUr
cjW2wWQudVEkwGMItOE6p8zYkqtqSekSRO+HsxbcD8M/xzgKO4JQvqS7a9zyjI55
QUhcHIttILJczFKIlgz0zQxNM4o13+XIXm5whWDgHXLbo5uwX0BUXBfnaLDG33Sl
n+3EEFz4jHaCJtGjqYpoHQtAYXeCRgHSciuPW3qg4uZ369j+grbK8jhS/DDrQAc/
IuoKY5kkXo2t5JduJ9KO/QZO/O+cjGPuA7oX4ARVM/WliFNK8lgDngluMEujFnp2
ds+gXGeS8GI080Mk6zMwwwKRIKsqHScC87oLID6cYq3osqGRDQdtp49Si6b7GfZP
N1AoBThex3r3KUPq7E8VV+7uaEm+Sj+F5gf5m9arXdP+DOmVZyS4plGT6NAWSl9p
Dyu8p85RCIsU2fViB2OE9IEnEY7X87jkkuzbU3Py69W/rfj/eEn+dwmiRcQGhunS
GOmOTMu3RmERfAOKhtQXBtWeiwyhCcF7MffxHe5RCgP7cmAGqX1qFhjZcBZRVAo/
AXXCsTJsW+0FqxIuhrGuIrR2fq64UGsrch5CQsm7lPu0CHSvMLG2EvB1sBrHM2sc
rg6hpNML31JNzVJlbBMRS1fjKUbk0L/H7r6HfdP8jYHuuZatI4dQcgbA5eCMKFUi
nllp3V/zM+GegKgogtxzrnEVACr3dUDLDq9nf/DhiCWi4w+tPbgIldqZzohDLbfY
J1RZqZlX7WVm14HAdx/VmXFsj1EFiFbT1dzOpZa1qGNYmIrYotSqAjKCw5zPiuvl
fGzyhjbLypVgPlVNkKx+6+ur/inVjAC0QzXpk2bP32ZgVc5jG69UCCMbHeKK6WYt
hHyNN9LO6aKGfwO9eBVa8DFxO8++x0udunOHT2IrP6A5cRNiR5t46zoew3gwCYh4
OcUUZICgck0wZqmcIlCkfrNO26uO2yl3j8sdXRdJzK9R+ZbAcuYxdxXAWlX6YLMt
FdObKCHj4h3gnbtfHmzxtNC77+WxuV5AXBEjsXcWCQoFZPAApmp0xwHX5B+j/dFi
UowkG/7A3yBSRYYjHMxlLGJGToO7HoLozXCMVh/inq42Td9317v1nXvUF97Kj+87
KrNA1UyNt9woppAhpCkfGhPQrvmd9E/r2+eSwwYYhReTDcrF/qIZhzee+dSqzpV0
ELCABajYIeLzTgUgTUE38DTyMRmjAEr2G2aR2cY5LnkdhSYGH45e5NHf7D2b7qO1
Yu25i0yxyrD+NTIGcmBkidiTt4BPGTpZhjanSGMbqGVnMt13RR32e4GBlyf7FTVX
PEOL3I4WmzD4DGIEMVmVz5Jh+i/AEG4eG7rlcIlq3fpxJf3OvKKZgC0iVC8SbIVw
JtohrMzjcBRqgGHm0+2XgjiLcMCam7wM2gZY82SkmhCNl4qSsH3Rce1BGEm7qXx1
2YNxCEqZvxYhR8BeOnUdNIKdxFk+PjhcQfPDvkeBluxA09/M6kY5lXmIEe0kp956
d0+7f78ToW645/P/dCsCkUlPzdI+XKYxdTkoT+iHnU+STZaX69Oke04MWzHWCxSR
MrGLBcregHYxCOs3M0kd3yngtGe8DDe8FoILVVRomhmnen7Zf83NHPrnftGlVQa/
4poFInlLeZgIajYacxkWab66281wlYk+9nqSV3m/t5ZmXT7BVobM/LJ2NB7LzXlC
2MSguZvL+pBTSIFrJ0tqpwm9ro47ieuAhEy8UmEA/OfdVh06eYDVTiqGFaQ+NsZi
8UgDYIQMScKDVaIN/7/6hYOXH85GFnAfjp1iueir4Eofg0r3kec1zW8lq8rTU+HF
aDSNyq3d3X9JhHZjFGtulVkYytPnAU19VT9+2DiE1IWgyKts4Hack6RUfbG9iuB7
9FN+/koWw+26FKwsewvTWjVUL60GBCoa0vYC7hunRoSTrSiiES+4ApVDfNRu7QOD
WQknBJClANLxckuGiDQ308CcZzAX/KOq4AasAzhnoeZjJ31dVfWNN4a+yJ+4ZNG/
+SwGrC/RU3rwC1omCWkFzV8Z996GHOhXE6ahCVo3f/glN+c9oK+yAauI84OGhOrp
AKdRox6SXgbS8XYO2bDqwgvHTSJhOySjK30tocepcZP5V1JK7IbHzf9YBAN5rocI
HXSfNo8SScIyX5ilfy8vLhhr6PWDvo2m6z9C/4iYJ+MHJrJUf/zyD9a5ch3Xg6sH
mcGgWFBKl5RSRcKT82hAjXKEH73TenmUTnxOphpItF514LyGpVfgz3TCyF3HpUu8
peduu3V8wpIFIKvOZQOzM7ORxuRY8Ux6J7gSURvg07L6T5wb7DkzRryJKTe9dXbS
Xe+U8q7a70Z1dko036NWukw8ZCCh6UUkIh71Zpj9j1QcuN9Wc2MGZii1XHFTwJg3
bHiFslxr7dqP7kKdg2ATnDN9a6AWu2fiFMGlKjLIkMg6seMoS5wg1H62O7m7whPt
MuOp3I84K5En973IcQePVikWMZBPMuh0+O14seTySwcn3BQeL18UFO1ELnVnE6X6
vOwJ/7359SUdqsSZmJkq1hY8zKmUrBVZvorgX9ASAmqjs1iYxC6bF5C/F177Mbw5
Jx8mWkvVwTo77VoZgHWZbpVlY4IuMdehU6eoDkzZl1fwIcKpVUto/6nwaWRLPBhX
RUoYnTtNgvSKH2Plwvz/wPmnXEV6OtD8NeSud8RbbR/4mFwwtIdyHKxQQVqByhTS
8NIQCobR3VuhSbYb0x9+k9Q8laJm7lPK4ZPC802pvwcQhp3c++mF3E9A4yYCNu9y
snlrhBC9IpvXtzgE+qGSA0QnxmKsxAlMtg20allQmV6v0C6HrN57Jzg/WPViUm6H
psLvPVSw3XYhbaPS37wQ9KLk/nTmAZmcjsv/UdqgdBsGMf79kIhnHM98M6oa2WhQ
QAUIXneym+dI+CjDfjevErlmePmQKj6balWmRNRgkGAFhbQU8p41dxJYPmM2slV6
DyJslEHplYBr0Y0aqOX7kkVxIQPAzydVV2DG97yMsbJqXVCuBjqV5gcsjWAH+18N
0CRqTMKJ16yVtLtcUjpFRO3+8/ylEA91Pdbj6e1yNTL+incmbhZhz3zaWSXYlKrA
hOVoWJDOj8loCync3b0wVbS4aRJAII1qm9bjT7HUoUQv4cn0fLrK1k1Wf4Sw96oB
/jcfEFJsJBxopu/R4ZmavljTKYX/DQs/pPHn1ztbErY7eqjGXRY6T5RfMtA30gBe
ozqKrOF1aGbQtGeMhMAM8mnac9fbA8qlMD0TjzcjR4Og328BLAYKciGiO142JB8Z
4ZPn7JPIRIzYCpFRyXy1iPuQ0MfkhsigUKHRZ+D2O6GV1UVLLTZF1rUjhUktGHEA
9TB6I+c6hSvUCuXsZQg73a+DgcgHi7ZPxrMPUQ135X0GXKBYHX+UJvo/iDj5T2jg
N6rq/k1WlUqGs39TiU61VIkaXt43ca1Ca3ewqGJdGvczznxqFnhYnHv2++c40it+
zL3oUM/PblfmIpXxQ+kcBO/RhTrICORwHITi6bB3yJp+CJSmaR8W5B36C9R1c+B0
p++FTE7a5wYsLUHUt52BzWJP6G42TaZNHykv7G4RTEaCatbX5Y/Q/Y0AdF+VHJ3f
RAzULF8ttN6KacsYrCnXBu+eiBsMpFbFCx8poTW2dbBSMErf5qiCaeKxsAIe+Pwn
LCSFLC0Z4/Z/cy6XS29lAKhiWxWhnuWC35oWS0sOdqgiGpJslwfMugpqYfthC+zA
5N2YRXcHkgiIEG0TOxfH54/O83pjKpyFnEm1xeU8546dX9mZmqzHkdF+W16B5RvZ
bk6tDgmx4NLp1kXYH+wXs2I7A3pCMAkVQdjDkyJ3bjz8R12fOU757/FWKshZM5XN
f/ADzcLCm3eMXV+UwROJmIsMkp6aiKCHpFbSfWEVcw36tCxJTYtpqbwrDPOdcNZO
6Zsp116u+YJamMMesOYtLUc2nNr1pgVlmB6jMqzRx9l3NojtV65S+DgwT46+ur4k
WbHwaM3LlJh434vbS+kBd+jIW8KdGuIVgBoSabumCfyYFDs00/+GHObDeQgykE6K
cHZL+X9qpmm8HMeTgnGf2c0JZIm4aGie71HFWIG3DfF/+dFaLLzDCElklm69swEM
UyWzvVf88X23PXXNFOWgp83+GntM+3wE8A43h0MgR9iAfoRvRHMS6+csFYC+qtjs
qgcFu9ilB6XMHlh7WTds2wjwtOSRvULFSKmHZflQgbYbmFceTVlnCVwgURZPZjnF
WntdrMxaLBelaY+DG2N2m+0vOZLEqwNFfe0EmhXaEOG0QXpR8EfH6tPupkz0+UmV
fsuePWw7LWffbPxbQXdosRefAKowm1b0BPt5KrEk3G8T8IKFb6O88SJ2GlL5rLhQ
YDkqJLsbpRANBN5fbUbEdymA7Ls0LL9q9NeJXGUjMNuMbvVO2fIZjS4QLGKe2E/G
hbrvfjC/KJMwGm8INtdjk+53GXNQA8/2AMjCfzQ8VN1T0r7z7VkUHUIo/1+op/Jy
iuLiUN25hyKYoE3D3eV5uDd5UZjaPEuwjPyUACKnlaOngUZKVgWe0PnquLk9CRH6
vrH5gsXvn1fPAjErl40N5E3xhcJrU6ofUwCGeFfsMth5PwtsrnWL0oXgi1FAbbnB
dj1MZRY3pRFLvjNXAvohAETF84NGZhCMqAavWLOxV0L5nCjc1GmDtqzd9QmhzQnd
M67DThfpViH2XHrFUTNa4YiuSSlfY+yRIqHS+WYpyXF7A9wrzzkte2Nu4SePhj/W
vvg+R99QTLYidB/sBKmVkiQC8ALqqV5lX4HgvjBk8qz1yhKQie2GeX04zLgOPqRx
EqBdMJG7r8TyqmmysdpOcWZtWAFY2o3NNScIluDzYKFTKCzOm7VVfWIt3Du9Ob67
slQT80m1EF5eR0DWRcEMLUTi957s3I4Y5IGBBueA+KcwkA8A6sR/ACrRcDLVUnjp
Dmm/Altqk3cUdUQPbVg6ZKEMKZ+fjis9eJKSg3WJlSQzEIwjndhBhI9RoiiiYoUA
Tjbn/8DTxFFTh943T8KrV9B5/CtDVBuUsTRqBFGim1hLfM02S9P95Dltez1HkNga
E5DpQOcHlxwyViDctjwHxeSLaUOSYjzLNXk4p5JtrzTjJfUkH45CL3KeFPlgeapO
M2q+gkK/DXXmmWRpjguaHM86WoKxVhO0OkhReMaU/fbSW9y0Tkfbv/tO90cHQWlW
CWSIpY8RwWgPT1OTrGB8XmHuvFeHuUqDBn1k5+IBI9vh/SJqjmc8eFRvF4+Qk50s
PCRkr+YGFbwCKPPm63CnhHS2pC+NSLOA5KGebgFveZdp/6YkGX2PBxBIYjr1GnS5
ycLGRXUE/qVJa3CwEsuJ4X8sktvSkZSpFHJGOEmtCwgbDm1F+2pIKh+Z60EprRAE
KX+leKLPDJy5KrCiZPsXmh8fiYAkw8ygDLI6l6MJyKDeLODo+4U0ilAN8HmlxzMk
YDZD6dcHpwfzOqaM4kICrz6H+en6VI8+BOgHS62d7CnvpzEs6PlzonJqXvs4Adyd
4peGDA08opvLE0Yzm2WZ0OGSNfIAbE+RFblvSudrSi2dOX7IFxIQrrFDZ3IvxyEb
w6yKO568jUOvvO5YNE4oat9ibbA1LMBqSTW+/jNcmX/8DYD0d5o6hdWOSMj6LLMv
/rHL4gTos23Ajd+e19aQu5zX9gE4A0wJpckOVsWP7PV6OtbHZbIxH5QFBVaFmqY1
xJQiLiaFcpEx7fWPGeHGi/W7zteRxMK8JWnmgyW5/lOaYs29dbytn41Z1cSCycDV
ZClF6pyj12+xmx4Cjr4ZmKhUWRaSOQlHd9vJu+nXWqLX/3eO46jOUPD2l7Y5XIYh
rBHR1JwMKbuKM97SBRXY5Eqz9DMGjet7zmDmpqyAIk3RTsNCj6EF0AQPEhp7MyXE
7Hhw9yaxiaD7uz9uVW4GiKY9QD0oM8d3x/tH7P7bViT52sPYST8qAPTniClGWVMs
tYJOtw51DHQdJD1Nt2UO+bvT7IWwxk2QMVZrGeAVF4coVf3pmVD4wlj7Cs+HPO3y
1Uc7eRVxLZLSDdRo9FSabfIi9+D8loA/Wl/6m5YcHJR2Y1W1M93spRqnIOY2Pc3L
9RJ4x2fzuRa9SkGerYMGpYHqtfFSo5L+3DkBF+NysKqc6Gw2B4DbNCJaDHIbxp08
Rq18olKZsAkrZLsmLc4aev/8gbCP9uU97LeWZIchPSR4SaUF/s559PuPe5HmfvQg
xxxvgxgbdvqqLkOHnApjn+z5U0Uoqmp2Fa/9dpl4JLT+CSWExiTRxKPUOtYyj7mW
0I8ELyO4pg6kkqzKanASee/ISWM+GuLgCOVVpbJuAsr+JhwTkj7HlolQCpXAqxof
G1rUXKR9rqsIcrYEgatMIbE/IE9+PvRgF1eE2XM7zpoyFNoHgrsguJO8bQXJyvKH
eGQFBw0Zbz16S0f/pCcGAw11QVtgMzWQnbWFen2QGw9a9JQMPXpTHVoDL6ZuB9J0
U6fPze1O3SPg548PnSzX652cTohro6KDhWTd6IhXdMNJwnYH9T+FCFEtc1bkKHer
y7ArWQV/T6jMAUSPiDRGzdEeLAfOCs0/oK9lb3QOO+i6vPb/KkWowH6ABNukq3L8
RIYgI0iCyCIp9W/H8y7Nhu6QIlGR2c4aI+JsNE3E6tkXCqoDIx/NiD6dQZgKGXDn
CgybOtZ7H8WdCmcgByt7DTi2/NN7L2L1H4757FOWtEMHIPDThGSzWlVbbiMjNKO5
v9W08qJWlhh7E/am7HTL4HOhEWrUDpSb/l0bPxQ0v98pyPjtRI1t+u3bl7FEwLuL
jsbtWD4jiHJ1HFX/kDt5d61OsHM6wbATEjGevBUHfmaUW++EVLAwYOtpfkV2YoHq
6H4WAniQOjEYVrbUec+/1/ij0ckjkwrruqhxj0TexUZipEovZJ5sdZapgDrlBOTs
/luk554aiVYQFW/QPBX0KzTZGjcuZ3ystUpF9dqPeBOFcq7iki7YGzkLJl3d4FuO
YtCCR9LLp0FfC/nArDSCePSiOG/gACAGApljl4yT9/IgoKfIolnzsGUhKFWiZZwL
tgDP4ibRwszSHw4qmalYeub+QN9/DT/jz7dQH/MnIhuez6G9tnB4qT+zqf67PG1s
/JYRz6F/EovkXh9/+UEPup+QeisfVY5nS/WO982RIJNIU2E1goHh/ZSjRH4KvuLm
1cKl/+kjHNFvwWeUzDR9k4wC/GstDE/pdxQdTJRSYALSiy3H1XrVNHTRjgr/BOGP
45SvC8x0pl9PCYmpebDIznheb7cTHzgZLutTZHTDo4UcB2fD7vIJsTL6EOXMlzTF
99+jmOCIUaq18DlAsEhhPuNW54gO7wTzgqgiG9TlnySAzUVtrwJzNh5J/n9A8csk
bfReuNPnhWhCYTjh9WYqLgy2jEJ3Lvfl5M3mDbth1EciSV7FjIhPuBVJCHNImbb0
PQPFKeV9faA0KkCGLtWE6jAlG+WPkxQbhOflA+cCpqhE90HgQsvpe+Gj+i2Y0ln2
LEBGmAWQU4TNyuTVPaZNcThk7bHf2I6rnbhn8TR96H2w+xezM+vBs3sQv3bDQLDu
3e7G3z46zE9x6zFaUKIiA4pJin33BMEvSIj1DY9Uy5ncJN8QSAaQ2xiI6oEFa6Px
XwI1azDdk7ZnWc12MwK+i46xyBwzpum7ZW+p6HuZIQtKgvOGX9D/XCuwwkzIZE4h
3jg2MlJllmDAxFmzwOCKKayrBmo/0PUqqPKPZ8fUmLLRa0nzZ+9l6hpCcyiBkPZL
0JAjANFPgM2PnsE4FZ2nOCafHZVFGAdZkcL1vUiRAVPrA3CYbabNuD1XIYDqphig
Qhrbx2djz2mxRIpeBR9O8sGGn+Lf9Ujpi2031eZcsSn4wgfKQcCm3DXDP7+SaD++
TT56PQHxq7BiIX+/vDCVnKBHhJvR5elv+enUBw5zxP7ugAALTOnKdK+THd4d5ggw
M7iltua+G85ApUWS2iw4JOV6MHqBmWEI5gfYkSD0I4qTLSb0nvJZLKGSX++FF9sg
`protect end_protected