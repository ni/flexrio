`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 8160 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eislOGByxcl/gRn8UziAa+H
mjgbsd36EQO5Ail/O6Xu+Xx/ROMSlvuBazdeHDaf8f7uGPI1OsOlJ4LCHbWXdH61
EQcjXMInU2MPkIPpfGuwQwIZ72KqhCFXayAyiSkffa957OVIZT0Nxo6pdguyvQrE
w+tzxTJqmp5OVkU6g+Hj+If5EkjJpW9GEnQ4fgaoNbg8LhEll0nEvwBwrzCeInKC
1LMuNLV+4LVFxNmWSFq75Oi/JRo2SGP0WY8A4djggmpwOJM2d36g0LR3j3eCIXSF
rm/IpRn9so0rR74Iu4lInkK+u4yYBihyCf0MOTt6mEdAr5JQYi3P9VivzxgXXJ1n
Pu0dcffoMutSA85FeEKHDVNYXjHKjm4/HdNbGCIRW9wflxmnzFqpRdoaMniT/5++
sZ9I51OwkKLt0gsymMpmWJY1m8dLE64cf+2jOGlOwAo/5LZXnhahkRuTFVysh3lf
JUcTrqOgysqz8Io9G+6/NjSykGvk0x9H5ScpNlvQiydVNFFQCuYuHSfOFARx/5wf
blTGxckT4yByTp7fMT0E0ZE922N7PuOR8V48j0jjH7Qlhmaz2JeNT4rugrMDT/de
RXqgIIpQ9X+D6tTmV+npBY5m1Uuw6/VTuhjeD2ueQxGMH6/Ak1Qn/Mv0MmP3lbHl
Qylj5fCs6n+SDT9uomZ7YEZocOajozcHup1EqzFq6X6MzyFe86uerGjPRGR/xnyh
66oQY1vfSIpg4Zel6MCDQ/ftBST68yUCHPhgqdGPTO4N9k3aiW+Q8qaft3VgXT4y
siM3WVkvDG99qySFQv0L9Q9xXNiV5sZXiDrxxasFsX/trJ7g3jqudz2wShYtHb3Y
WIjYDUZRESmyl5JUk6MlMW+IZIc95IyMkRy6Rg3QxRSMi/+MKs8fBHSTnW0SOW/W
Jf2tk7WFr/bpQzjx6im7lL0Gmnzh3b6dWQn8VsRFKLah5rZAoLLYORmZICFDXslA
gIAbIZuViO34Up6j1vcw7G+U0385ImrNSgWkw9JuXqU41xPbXi349h5VgwElOcPw
LYp8C7Z4f3D7uuTYazPXMjOxZ9KI3Ii+ZUEgg2zVjQzQW4EVV0EIj36GtRk6xKIa
rMwh+MDsRAfDarlxx+lZvzAK33R5wL5AG/2G09t54dqHLJfJzqENjOCeD32o/MIc
uSjagjwIhudELOPLGE2f6vYaqi8FyHTvjdwXz21p4xd0HiHQEnUAGfhwmSAt6cG5
fLBA2MJ2cU6Q3/X/xeNErBi4vbesjqPvqPkx5TxKkL5k3xhImpH0uHHsHP8/gJ3+
qWgeawW2E2NSPzlav86yBW2h1Wi0q8Mzg45N2KGyfeKgT7xl102dOnrWZ5f74C1W
OYjoMmaljx4x/PKAEPOsRLtGbOihoU0qOxzAomoh048yIlNIGWCK315j9sRSspxw
lFWUt2kL4R+DkDYwnMW2vqxK5q/Ifr8o+OJjJBvG9SQosetnDj/c2ZwaHvA/HFam
Rih01icTlaTyXqM+zpxUoTeMUQWQk52s9scI0sa0I+JDku+xRpzS1CCDUlERMwq8
PFNqJzzwv2xPwFbOjaVSglJh97JR5UAGuVrHUZprPq1+2BnuW7gBfMc71N082ybN
vpXKSUKR8CH/2m3T/9JUHIG68G4lF6meJo8sslpGtrivy1m6f/WKRxYw0Qvb+PeH
JzEzLHJFp9tpIrrcMjfZObqs6J1H+kfO4KNTnT+/RBOmi55UJXtgIbHAVa5aLLZT
AME21PJtqANH3DBE16gWeJyAkaQyjznrEzqTeMh+YqHeFaQF5pZpYJSo8H02ZiXY
Wj+M/nleRf1x+dST4AiVW661T2IJ8XCffYry11Kk/1vbuqWVqKMsANSHw3Rew8pJ
j19aiM7KxUfEK6IYqC2RRlrtMEvOVJU3O7mkNkMCwslnEHLzAwb/Ck0fkBEPChNj
ptvL9XeJzC55oGTjNo3XbHCGJ2/Cj/3TrHBlf49r9uSs3kmb24HZuCTNeod6EUYc
sYTroM/V70OD4iQDtoPth+A0+899u5lD6ohc2LT7o3V7x3h6O2fVuPk859o3lFMK
6K0V3xfR9Aah8zL1r4A9XUDo74FK1zZ4N8ClSzlTa9esCYrBJ31N56HyNbuy9YCw
Ozme2UROv9mermxcmO08RAqEA3VmgZcvLnne4mnOp9rd2SYprN3qaw3cggCidObV
uAMmm0IikooaNMIetyMRGeIAyI7++K/ndhcxbOKdTuYtVHpvmUZlVEAMP7RjiINj
33FCs7AdTIlE6gRlKHUDWETqBGXA9SiH9pc+KczKdrpnl+PS/o2UJJOf6GqhT5c3
nWipCcm3dvZ3+qeyG24yPCJv8ozliPUoUxXW7eVLFxSuhNb+aqOfXlApuGVELnm/
WfwjHOeaVxR4rkw0dY6JTcvR0i8+ysM1kk5bbjjh/YUwTGU813HoPav/cEGC1HeM
+gxdoNLr0/MlYK/dTEV/FeKjEVOhYfhSslT83iY/6/w91/zmioehHPK34cN1FXxL
mxSBEj68ugFZAmLqrNZzmUEJCWOzGnOLLDrQx7J9a3+oajMiJXCfwWoKUutfp/Iy
rG/AtETT6poe1vLyOw3K2oObbL6NpwugcfY5Iqxj5Fz5vDp5Ho1vZBzDgUsisKdK
hMa+Gj7Ex/MDhmMdKDd/oc1BIozaUbg2EXuGAVC8AQeUmt0zjiI5SVYIO0zy1V03
D+SovD44hX2WxK5tidrSR6e1vGVdfMoUQuFS9teq4fXmX0HTafsBGTyK9gGLX8qy
700P+A+xab9jldvPpx3d6DcTUKwPkDom9CGR4B0nPykviWTHN+mPLmBhsyQZW/R1
c71H6GE/Tf0JC8KzeF3rRetb+FDmFnIhjGlzbaXAgaE3BoF9NgYzP3GEFbyTEmZo
z8+kkjNuB/ZUO+UYhKCPESRrRM+DlxNm7fhoe+kOTul6TphV+aiaaptKqYkfxRh9
b2ACKiehzDRiij6rm6pCT2YsE0syc+ZuRjEa0YBMMAQUye2674YwRGgjm0urPrrL
GaHCqHh8miLdrhxssVSeM//QF+Wp0a6whWxQsyQ9idg99fbrlGl/kqQCLWBTJuYi
bPQVgWDWg2Bv0aRqAujcYpK+7Uh6GuPNn/lDa8BUeQpIXPJYjmqRcmEwL9Eb1P/6
PDZfL7L5rXWGdwDgRBSVc2UuzqHxlLHXPgEO3joFB2PB2J2ojZuwrlxKWUqGZu+a
+DZrPQrjkOewWFurm1zDswa4wxDg/cHMYL1ImHdZPAtAQrmMRTK2Ylv0UwP534QA
f6GzG/nui95XgR/6hPXLA0Q+2e/sCLgmay7DvuWRPELt4oc8N7qpUASLFLcmwqES
HhaNo3X80vFq1lNCY5sMVZRz2zSFimUo/3qp0sK4uvUsc3LKeCxukrjGmTgPFwh0
sQ6B6h/nQqipYu3NTxAVvMJXvqOQbiB3n3ns7Q9hvwE71IVqyvgh9Y2xF5MN2r6t
rJFWVzBgXi8IzYKqLi1LgaygCJuFTlCu8nBohw9s/UfeGr1djKMob9gnIaeoHRyl
lQ6IgHEzQ/7tu8Eas1MGg9FHxddauOTA9feXtDQ2KxQIWoahDbdTuKB1WU1pQqV9
sWnpcsHdmd4h309PA89mTIMTGKFvIzwNqEAdyWy/A1UeV8f8aJWlhpoq+hO+hVW3
wZA5RwalZfe4CDxo5zsiGshMFMvOW6GzZy73M5PR6ZOP4gEK3n2/aJVIUs8VXuUa
23TFYap0M0pR7H6LpqwTTnsCoOdVAtVPrlws0roNlwiCskDPZs1YyX3lJb5uupb2
BUpaMKkHdCoXVYeJwQQEmuL2W5riuQ4dZZA/gZHZulqcdbJEvmeiuOp0q7YKG6rU
9kHQKFCJZvC8x5hW20cVHuQweX5trJjP0u0IUCJoBvWzgMqtnv66R45SpVDS1wkh
miFqSXGwvjk6cqH+I12Z16YP4GprOmTaS+uFfllE4lsGX/3npeI1Qdt/Z4+KohAg
mRo41Nfo6p322nGvQa6koPdnHLn7x8IZTIEf6ChPqOBNd1qmCo3ByO/bjGO5trCa
fbWrrUqIeyE3+ZwHTLvq0610Ug4of9ePPR1GMxkgnbD97XO1Lb2mXM+I5dbca2PS
73TFgTDpyZOhX/slr83aB3tdK4YsBubbgIuAefbH5HyKz+/2mdgre+M23e2KqMyX
EFvbMmsO1waJCqUZEPEbkdA3fOj1rrJhVLW5dAWnp/91rYA3OfQ9NDG8fEArYXBm
g2RbGbtDEptgIulKAwVzOD+fgXG7MCzQPv5np+SMcdLSoTm4igxZdD9UF3Ax7Liy
tkY1Qs5KQIYwA3g5H5wstsTTD83Q5ElTC7/ZD5eatxdrLYH2CtXAgp6NilV86UDW
w70wNnOkeEu5p9mwoT9kea2AnV5d+SIngbNBCZo4a3A2FeQ2y7lvAuCzUHDuP6pF
nkkhzSJr1lnFemoBMnUlPDPpqRBlYd8G/AC7Roza/4nofhSZWDuzrwLeQu3li6hi
j6f6cdwhnuLnH1+jqNZ60QmX+gR8OFQKunQ7921NmElIoR3uslNtk6UuiL6R5hFo
+vemWdeHVBIEghYw9kznYOO0H8Pk6P0x9U68Bf6MmsXWqpaehNSOBV6gF5xlzYcw
fFLfGR0PCGeU5Du3kn1eN1/Ikl3VyjisTGHUVUZ6Gu1i3UGMWtORYB7KXXymRBWy
aC/44NDYFioBfk6UI5pzdK/p7ahM0UeIuPYjfdqmLNbyakZ8z0h7s+27E2MMyeey
oz69LUI09AdZb+VhffXjc4b1hdl2bc4gWVaa6P+lTXjFh77ufTdl0ZkU+fa//Bor
Op6+xD6VriGPdlTOc9+g+sgUThOmx4j3EYgqV3VxLKt/pqs/qp71bmbnfFM+d4Am
Ht69YUUXrEiydRgU3H/NuexnHuP+x+a7Wj7q7BRM31qwY9khZskxEmNdxoN903WV
AeEoSgWCg+SL/jHkMkQCOoiMbbl6l7SkbznioFmRV9VybmUxxkie8AAtiPoXyyoj
yMVCCiSkgAoMH7+fbod4wTpq0+kWi/zemCoqa6xbY8cM1KaL8wy0duAsUsXuXO0r
ShWWdj4AhR6TxGZPvkLV2EZXZNZjGSCtBw7U1zRXlK8zQjIDISojlrlLa86dDY42
jr+F5lM1eRhC7jIMt7U5tbnWdpgj3NbnUDxOp9mRSfri9Kgu0g83eorxDVHRbaRS
79Os7RnAw7Kl/IGD2wN0vbh9NabhW6lZF6sCBZSHnYk5/mLURJl0WofTmh/jxmqz
zBid4rHgz/OqZxv/qPsv4gkJOTPKGXFNb9WgFkMMGY5CFGHQjE5EvqzG1lJnI0cW
s0JdIWiyWQWFhHZfPlPuhV9qC+WTTy0bF1tOtwNkb7dD2/AZhVN2wDgyg62IFGJ+
4qmwzAaRM4MimpGiln3tKtFZ1CZL2RATTtiJTgV94NKMrvYmTLH+a1Wr4NLc1Iwo
HMcM4cvVkxZSrZVm/FSfUJ61MeXCn4GOecRQgqHT6M7Cjk6tohvYDkzzjqMkZhPD
V4S1Li7t3xoj/owOIUH1A8rqsRJEV0sQrTf3xl5BdPLcZpzL9IYMOomJpbZsOc/V
O9UAhNpc0pD7UpjyrYqbvpJ9y+w6weX5cryldCT7//L07xnWUFUwV5EUaTgDOKOz
29ZyEoUvXSSphFMOhg98Hx9aTo7VsfnNlTjx2x+wcvqIV5VIV0wpGeyN4lIDCwT8
hHGDdPP9Tlca9WE7v8fWjhO+oVPjj5jILhjTZP4kcSKlDWi9kVl0FxNEAMBBsiD6
kv0MogjQYMS7fgu4xatM9tlq0d/bpGys7jb59FmACg74f7es8TAOWyjs9abOYex8
pnK0IX/SzV3aa0n/u5WCUo3QW1VBVZ4G71czwyKykzDN/eBWvAInYs1GepppnEkz
AUBROC5YoS8sZHVVs3LbOZvdg8v8oXVB3fGzw5OGu54+C1dremdFJVWsw9JioimF
O0C9vu0dQEVpof/ZytjRZIFCzW0uN96Hu/Tz2O8BPzHN1A2hTW0xBF1tYKbWVo8g
cspYdAWNoELHSL5jDV/rdad5FEZtIoJp1bUu+64QX4Bu3giDxfjduzcCObc75WlA
J0WCIE0lqrvdmvhg0j7cO/iU2wo+yTv+Ei476bjIiBcU8dI9GKWy/ScC9+Cdd/kF
p7gN778R5t+iQj4lKsiYDv4nOAVW1hbZ0gnRwTiWFXJ+p3Zor0OiaQcS97rY/q4F
FZjjQWQaIZVNSmZPwH/FchgtfNPDp3mO9cAad/bvDDIDI6qxft/C491uXkuKE7JY
P2pv7zkq3mgcXSI3DWUYRGhXAHL4vMJ/0bXgdoKCqThvnXGBTjUcDV3rOlfcJPFA
31eBBvQw8Vuopqqlwqs7IkLxoQRcrD28RwHjwM9lPNsGaSuyNJRHU5GHojQAU5Hl
/EdH0rxI5+J3I4NZ5F37FPRGmDcf6j/9cRbBdcCevJFiw3EC81P4cw6izFAaoWEJ
UjPJUSwB23lHOCeW0KQhbUz/cc8KksJuYkaz504LgVlg2pX3dGgXPtGmIg+fwuCH
KOyuF9InPZZvsljC64g+kaM5MOi/4eWWP3by0qdupNpRTt8Em+sHcqqHSVlskQ45
Uo1PW2VM2j1laU+qSq4ctjMP09dtYy8h0Pvh8P3mfs180HHour64RTkZ7fCbS3TN
bSaz09nZ52+Gw2k4evPiG2zbGr6HlQCNyAos+WReXKzh0BHizmWZ1007L7mVkWuG
J4atxyzOHPjhgGS3LNr2kE/tmsSa8IXC/J+rRSUwWv8AiWj7Qob426/u2alZD737
ue7fX+n6mC1mjSnCqSQjq0KWaO+iSbHvz8FniaFzh2+/6/kjgMoY75co3sM50fpZ
onIJMxNhg+akncaU9riWSL7gWPC1Tn2P1elJOaf7Y7uy/uLgUGcWvEtDv2WeyC4U
Q6TRmtwMAz2J7DC/+zDEdLWEdw51+bWl0rJk1spGiX2U0dVgadwlqMnslWK+pgJ1
IQ+BGFXnchDukXT6HHwJsLiZUjQcPm7UJQenFS+JDDEXfIVojVbT37e+BLoJJTi1
BpAbG/oaSL08gIzUozw9fJCLHx5WI0+uEQy312qCJyIVev0/I04A+bYalAhKzvK+
6C8Pq5HntH8KlKBDY4HtDtK3XMr0VbUh9F2OdZ2cREk7iOHcY5FipdkeAVZck0vO
pxjhaBPdeZswuQj526BH9X3D+FCuEtzTz1tgE5/CMrTryuZ5BJbZ88hdEg8ArEkg
O8utQYrb2+Bi0jr+uZL6WuchBjJ3YvjEZEB07uBxJqHiqWYbdzqWGvtVcO3aoSza
rJivR5pMlR28uTwOSClIUJntAQIkdgaOakw/xmjUB9biwZdm+udpvUNI0yWp379/
XdEXZp9C1sGtS3qpXIEUB6eBoYPwaaAXtYCcx/x3m9Xgqon+iW6jJxz2rcRSQXeR
KW0jK+uOFvrPbIn9Mg+Aatc+85P2cCNWHjtMlIvUhi79wBs5LYbTo23/4cbi/iWD
C10i0rhiReZfnD5OIirRo4XmmoVbwb1Enl+m3XM80LMC6wOvY03ZURvxCTYC18l/
qIptuYpMSlGzKZ71J4SRTxe466gM3ihI06HeYOCyRB73afFLzjwz8FA/JAl9UGjm
+2wIB39YH4pT4hmRBYVdvPsKrgED3YmcrfahETVZMkOH5eXKqJEfdHRkNAMHIpP6
w+JT8VWYiOjtdLI07Hn9B3d+ZJZjIR5n5F/Mtixj7zvd1RAwVjidkm8bzE9hCJP6
jAvujmpsynotVW4n8FCH4/NtjAVBBdWdF8RqJLqk4Cj+X+KJOuCQUYsEuQ1KN+Q+
6yHWjXtAvqUgUmmm/5DdEN+fmhPQNECIVQWgrV0gSh8Z0zXvzZJLRWQy8lbw81fv
qERb5o681TidFIdHBjZnCAMqJm2EGPPJWRMWMBMt0EO9uipMj3uMqsPo3OBR5ZoC
vurTwKkomeR+0iOX83J1VrKn4yqqJIr/0Wu4PlSZ4tf6fUmeWntgZiuTiWPUncmq
qWM8jnV1eKi3Ao9lGaEc09G7vEm7HA7R5EiUo2lEhqkpuzVCG/RUJnpy2PS5tQi6
4VRX5LEgtPvGyGMepPyXsCpU+8bJZScx7tzeAaKs7WUNqQ3miWUqQZ6TErrNNUoT
dq+fl3Yd0jo/cyPsPLYy7GKtygru56QxWiiGJbhXwUZmX9pwoXIo1wRDDYBEWSIb
XGZRp1SwCeetQH07YIdjoJpyqcI9HQMPpNOXYcvgBjQibwKENDLX7iKeuxG0sACg
eiNcsqVSS5D4bbeshZoluWU9t7gGfofS5ri1SErKVj1q1U7FjQ1ueliXOM9Jk1vr
y3eMxn/DbUlODulXoCVlYvRJP4fqj+x7osazsfGLszt6vMqavNt12s0X3X4qFYGD
OfQe0fFbvsF3QhQ0nhLhSnsN/RofKG4Oz/paJiqdBdWePai7cN6fjOfscmulptW/
h5jV6RNrAd627ZFww7197IYDCBhIg7PRXObmn/iNG5yjdoOrq0c1dlzqnA4YVJS9
1ZoCPFwAkIutatvMq0RngWujKKEQiDKFI+JVIGSO2oA4cPspm6sdNhU6lkLyvhow
4J/oEVq0chp0PrybI9RgKDAGmn5UhShCLIVWHv2deiPhLCppJCFfp1b1RrQ8ey0l
eXx35OsUyINVcM9hIo9JQj+8aAlDB1utZvaL0AVgrDK3GAtVvcoDaU7YLRBIpc/t
ZCelrzbWiZSdZHuhc21TGDIN+ENtc8qZTQfiI+58VPpDO2s3bkK+dKqPC6/e1/CB
B6wdhwkg7AmfZwLvzJaIumlFsjkFx634nxk1JXQBbxoQIN/62rbZlKJZg2xUWGhS
UimovTuab+2CIYedyjuiTpP6CmvRxyAH6bU9+aIbNirFMNDCSfsRLsBDMpsFAR8p
+KcpzdSTvTsZjz1ZS7DWBHICMHesxTCDL5/dzZZ+F8mUiaZeHBwY0+12zM9rbFcq
pS+ifH9sjbznH1YWVUNN80+njYP1yn5DtrkA2OtYTMPbtudJY92VYbZbgsfBCcKC
nY8Oy6LBXFK2CR67l5S59V8cQToY372f+34ciuViLrThxPZ+jH6HnJDbF+qUvRYQ
iIXcCv2KNBgEUPgxVORCIL8P56vWA2h187ZvDLAN7Xo9XhJ6B9Oppf4iUpG7xvFp
apE2TDZwa73M2Pdlix/QH6Z7pXThSF/NU7WtUbKEgSCs08T5jd4QbXgUqqwIQe/W
UKqeDO/MWt1kpQudiEw+kcjasjk8L1jgOpyU+/WY1vsxQupgusacUlbCBF4sFBG1
DjLGQyv+93TRGD2ILo9VzxKEuH6hH0166KcEYXEw61NOhUeVVDwzTIgFJsvW/q+f
VPuzqRq0rCayqceqcUp90CKhi6h+Cl1xsX6mgikaEqRTw23HljBWV/708hVnx/au
qoFHhpovS4s8eVzLBNs+JaXQmcliBg6bMStOAEiqFJ/9YjqC+jgXXDX/ViCIF6FF
lpQcCrTzDN0UUa5gL0pXaJV1RP0e8lQw0mTw/1ZnwWYA5Jh8PfQLd/bh+6AFP3nk
kUgld33utJWSXziJfpjpgbjuriLyLDcDnlusSeBLvsSCyRkZW+fhm09hvdKSmdm8
eMFMkBwT+fTJdsGi3D7b/aviAnYqARM1sRiBuGCf+JXQGYuPCDOYptq1PBejhNq7
fhaRkkLzwPwA9RZHxU4ikVNFMLc8A4QCZwC4zo1ZjQU1wFpsQCO/4FQIimZRN5+p
PTFbp1Vx5gC9runGiUeaCesQBcpyBUSwRVQD4wIzaTnMwwlobVt5G2tZva5XSovz
K3Z6Q0Oyf1ZmWblJ+Pamo0oTQG8qFqvBCKhBFIhYbVmkwI5yIWpp7zI8hYHfkwks
gdtZjlfqzlz7MpzjOKpVruInIiv37U5MK6jh6OYCyyF6yzP4P5xb2WD3Y+1XjPAE
tpvWWbx1HToq00jV8EPo3lsVRa2Y8Rrk1XBokEURPtyNKo121yjN6HXXpxA1GKCt
luUDFHKIphIrY76oh9iHoSUzCsIoWbsg9yrDFJiHFpfxGKu62Ph5AQpP1UW0USmI
pUDTN9AOxqNFVJXbvoKWvb6rLe+sAAcZfvvb9PCSeDBiFQBhdmkkw1ornAye/u6m
APMI8Z0VZxZsHj9erXU2lvNsEzmKzzAEk2LfacXfF+yqhnk7AfgkKu00aFd7rpDu
k00feKMHNepThqMabdrabtAXIGBTnH8lQyUjKjFD7IZNDeQAxXoP1kkX9a9Ytur4
bm7rUPXdhZQzxMp3OCmbTgiH4RAMWMu9S5AgeMr17Lhkqcy25BuW0zr/ZTLUXA7p
w25yxlp4rgKVK2xPhcpIpDDSRfO0S+Dg8rxXIFpeRKAhf5Swrebx/2kvDqF12VaD
QdMmC1K6WauRPcsRXL7IPIJ0v/hZYCqJETC3dvDNpPxzHh92UzrfkZn1xHRI8mNZ
22vpxo6xhwqqfAg7z6msigep/YkHrYQCtPf90jv045sJU+FmC0N+uJrhqhuDqCTu
GSEfFW4zOFdHxx3ALI+Kh/0YIb+g/eBhVo52jhb3tzc6d4POEAKwtEOsKoYJSeAH
J++XZwCRhK3MtIvfffW/vfe66rI/N0zlfZLdbDfgPWewDFKvksvE+OjLfXFVgqL6
eOWakEcEPnplhsQsCgkcJUB7nshqtNRCVwnv5BHGEFE0UKKRIWvFKenazTbHuoVr
WKHafz+3/o87ZWId0TFGxfZoUJ+yn3tjkAjYzu/XfYQAJG9EMGKr6LEulHG4qpwK
`protect end_protected