`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 13312 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
KKcya8NExyVaoCvctjWPKZxVehQchGcFvWDRL2K7qhawTDplTNmZ7s4kaERRji4Y
E11j8C3aMv7FUMnbBlWmbdCeLDu1jm1jdpdGUenxlHLorym7whiYlRAbp7eJKkqn
5i2dbsP1yrq8F9Hq8DyuzvXZ3ayRPHdijarzoFEIiq/8kFovi+HUUK1mTtx6+mPG
8OOzNVBdF5/fINVnHkrTmAX620khb5NtAQMqfqNKoU4DlQnW6X+3dm6x7sHuiko3
37UKO4Ndeh9wQX9ZF81lVmGP9FMfuDCOmtMAFkniyX05QLQwjuh0fbU77F98JQBx
/tlPU3Cxe2U1RVtUsxVidF24dT+rhsoOH6QmGtd5zLbmLUnnqJc0kjxEJ43VWzPU
ojs9iJB4pwTRNfTbMEL02SbmTmb/8FtJOlb0uxUhh4TYOC+0c7xV4QpouuF8LB4w
B+Fg54/74tnBYxOXUeAKNmIIDqKdLNN3Gj1kUdFqNFNhZJVrF3va7FIFujI6GMS5
TI1stecREqm+jnGH9oDWFNBdxjfbXbohQ0f7MLRzZHf9xGjB2AeSIc5vYMd1Vr7C
uDIz/qODMsqUdkG5g1hsSaaRyBABRYx/MTkqrLOdMfyo0mTxdzE9y+Jm3xC/qaNt
zONsoduiy+s7i8N9cA9sWydZfqrY0Ttp9lIleSRK0vxPuQbXdF9TQiAsa/aTf2H5
K+b+20JymP60d/8HxCKM/R1bv6REELtpZwLKluDRIkURIuw6POHO7aGABzEzA7Xf
+6qKYwcZXx9FJh7Wl7XCTtEnE2pwfBQuIrcPe0A1bE9rB5W78223N9Q/yw6NMZex
bz7Ux85EYIcR18c/JwwQDDAvzMPoEkLhtSVZ2dZ+E6k6IqdPwCL/x+Bmz9jXwD4q
XA8VGWjCaDY7p3p7YlTteHXb44IDujtUj/tWYNFZEqTDja9bahwSwVOf6FCCRJ/q
Jmb5mbG3Up8r5o9U+GIq7BPQlfdR/N/ybNQRetiFxwUa6AD9j68rznai+yW11v3H
UvpL8jIgJy3C5AIbcwDcvCe0iDXJ9xQx3FxlQ9IiOTMtgVOiCx8xDH0qtDGmIZdY
8ToHW7aF5dKN4Hu9JGY4rMepJUXn6LRSg++t/4aGVFWYpz0WeM5E7vCljBo0Ldph
uUbOz+RgoQzMgCFcW1sS9z1SbrQ0Vj+PVxeA6Oj6X8Hv2WMF/Vh12f/K9odVs93L
3C241nVQGbjbhNXswdsIMocPFuPo2/P352rbWsY1nOH7rCmGxWAUSu+opu8LIfu8
NGo3IKZL6fRPqz1bJjXyZtl3gXiA5D0YpbvNsrtewAvfbeNLg0ez8rXTO4sApZ05
b4s6cGOYh7TQIJ2t+18Vub0oa4NO1W4jaoyP0VP5ajYgcHuCNyIIUvh7wg/YJKAi
mzO70muFfe+KZ0Ggj+4zLJfivx0t+eM1GfyBQB3X+UqwG2rE245UFZh4pgoOrUbF
a0YO18AICBC43kSPI74yVfAVgTZEn2PWwJS4C+64cpfvF+nO76NLnWYMN1d2t2ow
ExUbu0rnTiW7je2VTJTCNgAxJ4d5PEXCswswip4xMN+wcOAWBcSs8ZdOsFsAr8vl
MJnupk4GhK+KL/nR24ULAhWZZrczCGbDUQry3hEk8xKelJu3DqVoCmayduV2H3cN
Ts451EouEKpXCnh/M6h0pClUaEol74e0AO00VpNv9Ux7dfsLBb9mpT3CWSwCCxdt
3aDX+NPYhn2gm46aSxgcwy3d7+QlKh2KVgwXIk0wf3OFrhs5RQ+G59AZ7YdB/L/j
m0+YoCm2boev7tHdfj6BYCeRMzZku6Pi3Rf110vPe1jBR1ct1v/gm6/V+Qx7bHtT
ugDzHzP4+bAlE0CTOs380bGw7bumkxp4vHwxdM05HpYgEjQnS/gBhZeidecGGpZJ
BO0ab+f5IVtO45v/nxgzxZCgbonF6SfibLvJG13961XkHte4NFugW3CBVZaNDvQ7
AR/nXnNS2I51f/r81HeJgQRIX8g51xbcXpvK8Kg61G5nBJM7Ia1iGJD4WKW7N775
m4zwql3qDbtoZEC8DmUUHpMtxZUnILU5JWDNUpqKii8suz0ZZTAfwFVJjIDBYYZs
2sCFrWNuqVtNcRTJHp5c7ZgG3c72HcbVHRho4WcdSGPdbmy7hyOilaiudN4S/d3P
dtDHIPF9yOX5wdzhvnlp20O3v0Ayty9ZSNujIMceY4QJIYLtJ7O0LQRWwA16weRV
JGaD7SSeRfYV3c0roLk4BaMSrTGNaiB6PxE+8NG6sIKEyTei0i24OQPYY8lPiqby
/gsoWVSkJ8Y0hMmdwTcXilH5gd5bTls9dEdRi/oB9DessHRnQfM1WTcrJp2hOYMO
K/G1FighLqaH4zp4pIynZqSY+ZAB9gIie5TbFj7lax/3zYaXDuM235wDWfDDt7wx
lbT/8zHWEdr5ZcB4te9/ibcvbOtg8apr0WXp/gn6JjFcxBs933wra4RQwQVNj2T1
ljys87yAz+RSjqqAn821MQzJKIvNzYXS1o5lw1Lo1MngKNNtO1qXLM8fTikhx+Fp
gC/7BVUE7wQM9YPh39ScJkH/+UPgpIYJ+FaYFL7s/LKFPWm6z1QcWGq61yX/VNBD
W29d0K0riXvUxjHrONYDWtcbh2c8PlrwxnTGkIa4VkCpvWpUzo1ByHLremul2Gi8
PmPN6ykGsNu4KUwca9lWSnkHty8CeiZGALfMwP7K2qiYMNn259AJimZk4uN7W/ii
d+fcLbf3bFEGecZzOvVUJciCq3cxzWViRa9CPpAR4vEuxKF35vq5D3WqDav6UOXc
/SRTWeU36PZE3UU3e/RPS0GIvmoMakjbNQu5u2o5CcN0BwwnIE92fiFa2htj7++J
4b+CdiFFiOzqcIDEPpRFK7Qo3sTD7lqzjo+XLn8O6a+4tSdvwgnF5KYs+JzCqsU+
vUKJ2XunQtXKP5VxYKvguZgIG4+hV5C2gjc5WnL4gZYndLQaOd7vc72IayXLf2Cs
Q2NuGEHWjdf2LkytcUbkmnSwzqXwRPBW9/oRz3E85qp8r/33XKK09sj2w1MzsPPR
8L65Gsldghk3R0JdBJ6ouuUMH6wyRfFLXG7AftTtFFv/G7njSL3sC5ZsivLW4ilS
QSUrdCfbYpESKzeU7mMdXpEKbOOYpHzNcUp5vrYKepMk9GpWUnqKH6Z3HkbylVga
19+u8e9SebyJYr/1lfuK3xc26ARf2ZEAc0fc0H+Ph508A0GHg3A6KM5rMUCjXdJt
ZSJDxl+zQFqNpjrqCtt69pdPDfvkeehZGLhLkjAx1x0MEwpIuqcsTc2iiphA4H/1
lFNcmvSBoG+X6S/Ad/MEyUrQ4Wb1NIHKhZ7NR7anbcgJ4LmL2vAk0jqUuIGmpchB
4Z1N5msycRsXthZH4wKuVEFKVwMog5O5br1IazKHeUAD5bNSrgV68fjoFwWRsIZb
AWIsY3r15ViDJT96XnT2jFYG8ANRZltamgzc7MjWhKZegndSNZ2yf4mtlBSs/XiS
nAn5kQ5J2XolQ6lUOe+yqoGjscbEG8g2BDgn/w6DmQcun87DL0R0CwUSiVRpTftf
J0DDEv0aIvG1vwkoJxD9G6WtediiQRBFGw6nn5c+JUmE9vdy53DZydAhhGzprOGX
6SNTMMV10V9dB2JibL40QeLWLe+GPzWQ4Qnb6DjesOxtI6Ww+Wfc6bDS0ZaVzJ3/
X0SAJ+4U/rSnnZskigq76Ju6Z4NazBp0nzVCzywd2OG/8Y2HIKy2aGCwwqhZV5El
vrYscrsEjkg069IbTqPyxY7knF78RPfkLMT925ia+GzBOfp1aHsVPV35PcN7IhLx
qndCdP1G/38P7Ke9uD5W5ercuqwONnICtgnbRnAaoFptbbFo57Z7GOVQZcpZwD6y
4crKmU5fgLS8APl0mjASaJt6dbmoTChvWDrYnV7ksYRuaWhYLu+doWTgke/glXYx
EOUVhtaX1XodE45kFusr38+myZvOcqd79Hrp1vhfMfByictIa4COLCukkQy1gUsw
qFcuefkIU8iRh9FtiKTtqg72MgUIzfQXYuMiX9hOlMaP+rlCp87KhGkWlFMsLFpQ
J3HhmAYXBhDrcb6xUZ/nsDf9LYhLngce2ZRTKvojQKDzJxLiBsmh9nbYjlndMXKB
SPXd1RHhDfyx91lOo0dYesFz4Zgf2vY5UbocEPU2SfaBSSi8m/WqkQMzP48VJyOX
OJMctniFGZUOiR4eRswgRX4Dn6H54cJpH9SOvhhDC5e03AUIpC3xA+ESZGII+7mS
hRnFyqQktAmdKUhmWhWsgprxKIysFKHfx6oQ4wFfUz1aBGkxYZ60UTKQ98s8Kyrg
hEFzWKdOEAou46ESztGU3emtyxg7uLt+nHskpfNNZheX3JSAZa52xVZ5pD6s3s8N
vslbQM2WHvzrV+yAmbxNLbXTFonDImf2rmYbOMmEgfybWRk3OVRWYYvaXuBiixg7
NkKK3h6b+HeKWF2Il4eFrR2oD41hyF/YSS1VrfjS16cKdK3vT1p1cptoqsELSv1e
fobQE5nwRUOdH6QSMbepKkE24pz+M4acacYRo/HVEvRLuYLp1s2NJwlHZyKVBgWC
YKWKEDvFEdXUqaKDCgQGXfgCYotAW72ED31x8GfoOc9iYbLC2MxLh3u+0S/pDZEN
Bz8/cJNgiDtdw0AJx+s7/dNF0syv1rSoxTA9Ks3/fyQwTDMUwyZrqMpREqxHXqak
8Y+REWmpB408s20mJnhxb+MH5/f/4vFGB3iMkgc5QcNYsh1obx4BBfygYtF8AbK1
rihmtQvhooU0TyDgI5EmeA138/igxZH+dXEBG8fOjR5yVgsKWAjlLtjxEkKKOxjO
r3jeSbB3khFPFzSZEB0Llipuma4/IULCtPeDBE5lMjnbXy/ur4Wx2NW56dZnJ7zW
xyJeK3xcuWugyfCkBrG0ZQ6UxRQXSP3UgcfVTmnoO/aF/5X5ErTOWDyCL0akxwHt
aCh5xOO8ydkChmeDc4+FK15mQ7aI+gbIM8VqpUpSkjEW3HjyQL/BRjwwyhw7cK/W
1wvsF8naERBzrzytUPCGt1bL4innz2AO8OnWkG1Ii93i2p8751DNqesEEj1VdlYr
B2bedEnoUHnM9f/ao0u6ViqWSKAamdLzTV1PC7Y25A9rM+eqy+7fM3mxJPvJI4ZI
TQ2ebgvmF4shsddSb79R2cwFJkAlS6qinxs5dx5L8ziQHV0X1MuUDoirUEHLaLhx
OWKsR/kRUwTwbqe688gNf4YJ/DZMKaqMKd35wu6Zxja5roU5IKa1eReNlSIavbj8
Hmt2r4FzUKFU2aOYGmGqwgxxm8KOCORTn2n2h4BZrz/G2p5Ta9YutQxv8lQTABbE
ssf+DCiuYcqhEUbT8/8zzJyuQUc87f6bOCo9ddWZzfDOauiz3lnL63a0me49P/j6
aUjzBdSVLz43V7N+H9I8IDOshsrdNGLz/L6/V9QgEPzEePIR9mkfw9mhGXjC3qKR
fsYg2l/JzOA5aWw54u3JOCqq/fDAidHiEOY/iV+tWc2YCQXIIJy2wc2YapnkfKhy
gO2sVAYor+vhsFK/uXHH+Q12OOt7sPNI2RCzT74UPcElqXIQe/nOjwrT6LJA545R
adl/vmyJwnkfL2NStNqQehh1f6sTcNXqO+5LS+nvpYOU/uZdEVPCj+46eBizQRyv
fUbIxbY8WvJzLPPG9QoafwwNQgRcUfTCN5bpFMlEPUjMKEU1V5j2AvM1Pu7OHtTM
HdbMpRR2C3LkrtOt5rU0DTKJmyqxNpYZ9tYgPxWeWZyTrhpZGKKFZYJrTmNcBRo4
cB0k+X3ZlWFPGDoCWOlejAu87XGOC0GWybAq8BjfXncIMz1GUa33afNdcOKfKn0A
95zPa5nmxaiYJRy3rjGD4rni1/iUgZo287cGvIWHasT9HpG6v171fs645ydxFMcU
7tUKF+qOJ6iCrGUk3J65KoECcCvpZ7fePNrSeG2t+9GLh2ajJSojqDEq0ZMFdTib
wAiNoXdkP2eTtHCRJLwjWGIWIhbvwVB3se4+GuaqK2v344bFnAwX/U+7lFRO7i09
Phw3b7a+8CPM8W0gdGYy3xMIwrxjgNa4CHeGk9w9wSHrnyzRtDphr93gELyroNNW
2SXBVkMBx7Q2Vz8PCFPNeka9FVoFGJ4Ndd9U/oIKVSWQEHjyVARQ6k8iUzNGRbCd
VBmT8CqkHmomwT4+11Vf9CcOAcp9RFKaPqqbSZh9X05KW4HvMlC+e2B768rduUAP
18gowTMB0WeHXzfLMWckpL3OrBFwSLx0htSN2li7DBAZ2AwMitEt+P1lobuNh159
mTVVatUJfYJ9wzJi0+uJHc7Xoc9gR/a6NrGct0AoRs47ukFa1Y4b4wmWub3S0my4
WE5z/bb+41H5G1xaF3vGIX44bha8rz2oEdlFFGJzxMi5uIsKAngTXqSoddzVi/Tt
Hb3Ubc6HTgDRCl0/ExZRbsoQQfYYMPUHw7Na5qlF6/qxzoK6AzrH5W+4pq0f89JK
AYpwK/wjrzVAj52HuyPndqgfWQYSCBWgPVc5Tot254VUrfBI28ASEuL2LspXkX+4
UC8ylBbyCFQ8q2mA2/pjk7t6wFRNkbmv4Q0qRqpingTmngh2C7bMbWQSjMPxSoIv
NMDJETfRcRgVPxiVdFyXVud/bBSzSF9hPIsYwKMaefTWzuRA2a4Gf4KRxSLqbum+
9ozJXqYXR6holqY4eRjzetCcEoot9ZmteIrFRPFtryvsXeli8cGLjNqP0WqHC/we
ETpCgbLpZorE64e9G5+bgT8BREX+ngXt4y+/sAaj6iezMhMh185Fu2uAJAV4khCV
hnq8yFkRnng3k9eosbsZ0tujxru6W9103+rfyt3orCCclKaSFjGY/fS8CnCMSssX
Vj9AhLVCqnYDHNFYTUiV6W20YjPubm0cL0SHgrtxQ4ws7Wg3aPAH666pYG7/VocQ
LHIzh5z7f3eGu5V43AUi/CUrqL0W8QgpJGIuLXcbSLKH/INOxLYaW3q7+iNy7gFZ
v4Bsj+/0RC5bkJ/gszyZRvwMwtJJaFYX+ISQPPNyOscsKPUcNqsn56MlQVM6b65Y
6T1/BWs6en2jlM+G3TpoxrXHfI59dJrhEIyViJf5nQ45ePG35xZzU34aUAc4C3gC
fZER+5r4wcPHtKA149Jfy5kAOi30lru8cSNVdK49jTL5Resab2/tUFv58hkS8Cm0
YkuM5MBSZaTaBXk4vbTQXyu6lyPtATW7ZtKLzMxf8mtZNoSb3K8eIzP8ND1vNQnA
qp82V4TBkMIuKxCWs8GaaN5l4ouzgjf6JkjKh15DRTFKpsyDHXY4hdmZgCpNL12n
I93Qh976NETPf9HXVJd20n2r04sovZ/y9odV+440JrdVfClMwpbk40fho+rAzL9X
sa2MUMl1a+F1gavsqhGbtJ2hXG6l94z1MYTWq/+y+enMAzAOGJikWPncyNeeTcMx
7URPv0incFwAZogDOSpGcrc9zQ72y+0CENjCuoddqhxCYbq/Fmo2dBUORYVeyDrG
w7DkJKcZ+m2ihnE6lIbI1AQtTn24DQVJL86ceGsfHpWYTqThft0xiDdyWPkjseds
E0EI8v2ZWIVCP8S7h/ehDX9X5POBvxhWB3yUibBvI4y4YlTLZxNSLBd/ZbF7hMOO
AwrbQgYQzehcpZQP/tHKNBA8Cqjc/0m+kVLfXRjU1Y4l6KbDZ6uwX5DXH2PrcZmN
HmvSrATdZ9/Ogr9LtdaSHPio7L8yNv0mokukspAxNoJ6dyDIudM+99kf7/93omi+
2qYp2iFyQJ8Etcq/ZAk7W+WT+5Yd6w2K6CRJi0dMiCucNUZWkLI5prEMhgb3hZ+U
ZlZbUfsmL+faTHvz9nliuf+3cgphPTEwevlNfQtKwZcC5zzFuej9xAS8hqo2fHwB
7PJ9PXfdaNkbveMuawK1mWWTiBIsfJVv0EEJw/0Q1lMdsWRITSip8U5LE7JVxmoZ
18/5qThbC1qeRQxKIJ9GJMXilVBKgrruKiafmGHmFMoQo8VS0+zNqLUnZsaMyIrA
u+fZuAg1vwNoqpi/ZA0aaeClhZHUgJ2xAMwpoOEpJW1tCqMvfHJ5AhWI+LAtWqw1
R4JYQadHxEyY7y0QaHyiP6a8Ew9LF8FZjcqDjcr6n2hOuEuWUfufBwGxqynOeEey
N3Qo3fajCPgYScWZYvG/mNzSTWQhXZ9Wr0PgQiDNyae/bulXC45ms2KvuKPTfWnm
bA4zVLNwFb3kjIGmjo6LmlWti9ePpOd9TJm+3u2G7qwGItfzlmEbqIFt3OvQxbqF
q0jojiiRakp2JtQEerEGkc8WEGJGB2dkH8lFXCkkH6YdJ/A761L/sbE3piyv/f5M
mcjw9Ds1oHTP90KwI5vSPfj/7oRso7R/f7zKXJSfyjwf08MMjuPaX9zKDYXZDeQ3
JNJJxRt69+DOXgdQo6nZAK64z9+ku3sQvEkp9rYTSHL9+rfUfWnJOA7yO/7i0+a4
JqsVpS1A8qfRx36Dt04MyApDNF8eu+OFDi9rELxHGESnTOYKJ9wVffqW5LOOOrIw
LFZaFDNrZGFjd4KfMEl415MfrZCLuLyIxd2PQfUVYKfR6hlyQFn6PnwGWHLDDPEG
eXnoSdwmtkhBs/Ouo6pC9kRyX4gAxkwFiVN9At/AYThJvVNTHoKvUq+9hvnkEM2J
qi5GF+PZeoRXg0HKSQ8HX4f8L5p5Lj94LPYKJO2nbyLSxWrv0JbhIf0kAZsPIei2
ZMdxNs0Sbb9PlPnvLxpXfqQ6tgS/d9C72hsNfgvJoJ2dRZq6Vxb8kTCfK3awwqlT
PS65dGpR3OAPt9tgYSVMZh5voRGW5tblyfoqCcB2N9+GUhFErtZTaihbNWiFB2wl
EnqvWm+PlipRXB1DOa2SBUEah5r51z4hxnhdSEWyhPGxzDs+RVXcjJOR1mb38Qwd
ydHf+i7tZHkTmUkosoZFdqEXeeuvfwGHGc7IGdOVTw0r4qp8iTHUVzBzUi8b9q3M
gyyRIGkcWRoCMQgqwIgesjVhSd89GWCT5GDqR1OnHVIKWmOVXjir4AfzqnieK/Q7
F9VtAG4uUOZv7Z61j8acWLTyxPJVX2Yo5vedq7v1jKEcvjFDTKuR/Rrr7i63HtEe
8QXeHAxqyjMjOTN5bNWsjY9qjjaHZoXwVAzu3V7xuYD0E8mM0L08/Hh68Yvsse0N
CbQc6u1R+5Y6tO+P9VwoXWJbqDHHuOnIH+rvDaUd4WmEFOY6CHNkQoDr9//Jy0WG
0zQxYUb0q4FGrUIh9aZxJ2NcNs6RTDE9/W62kky5RcphyBn0yJ1rGBmp1lykNfsF
2wCIUrtO4UiIu3oJEPv/4tmxvWmqJY8K0HgZDXTkgp5IZbkQnpuxM0ZiVdwshSv2
mSu7P2JcWMUx0k3p4eBuUK5Af0cDD6zbApRnkZqepx3BI4sZIzUODedkysCWHxJ3
QlIMe7KHKtGyIDRG6/cSltiO3HiSVo4JHGSmK6FJPuyoJQaZTw55vX2tMY+rSiN1
IdaWjI+w/wSKPYMW4FwDC16ygubOlU8R59r7fa4d433/OH4n5M0dw0J7nhyvhGo/
pfuIY6d1VDdPz9H1qnnnDv5vLMAj2kzow6qFQpu+E73XXl7BYq4d6JjS4u/d/DS+
2txvWL1rH6/hs+vlMclvD80THRKPTivrOdeUqujckFidTZOLdfDCS+ayAaegAa7C
9O8Jj1zM4in+nPpnP0C5MaqBBpYbK7WMSP7PfYm/ZIpWYQjIRmU97Fhr1siLGI7v
GpYqS+Er/ptKVGkF9vxhCgIFn++UwcCIv7E4ijm9RkXELkI6Rl0IJ32/4IUVzOAv
tCPiY0/C1bpiA3vuA1VaymjZWTpFoiNeGtSuDjKc38wTySRlnPjqlOq8jEnxWiQs
68pdx6nIYlB9wFRJ1TfOSYwRajzBeaRTGKZ4fIpPNeI2qtpQ5k/Jaw9F3266ILIW
XVBIUaXVjYrgR2WOYm9D6jVvdAuc5ASE6BVaVX3Rj68ArFsNXe5++06srLsQeLkk
FpnFTWtBjvpYtPAn1xm2sYICk8u33PCpo5XhsfDn1oxEDISSQb/hr2ekyZ7TPhnZ
Kvj3hDInGq74ZP2DRBXxccNp4+IyTPnmX0TtXQwW/RHjd4WsbRS8xxVheIMyloh+
XPHU5Je+lgTGnJTKnU93D3EoMIT2gA6l8bODrQb0Kra59luGzJWV5ZSmeLHcvAYE
dtmCXA7RYaCWYSbq4HFP+KWjmvprVj7wlULerBoBaqU0UTMsPBgiX4oaGZ7nC75D
3AaigwIheTPYl8sVo8ixxzOd76PpA22Q8g5sr6OGELKUweRu1wSGRl029PLqMkRz
t1OIsRUOh1CVkkVYIylUP9Os/Ac4Z7ZdBovXerWk/8mnJkT26vjPRNofmoOaSuA5
DvAojPv94abAD2tXuU8N7rXrUceTy6QT5DwSzfD8w4n0KBDdnMI5kwyMneMqhaWw
M80KBD80kiMYsRhD+SsNR2zQH81X9C43gTkL7TTDF0nmap+kyq9Ar8ktuWetXaRH
yMmERu02yZP67VgUgTgvg2ap1MLlfBkKejEeMTw8yekW01liyfTlpWXsCjIrRDYk
PLivzkpHbxQoK7HL9B1U0NAhBjWIlO1dISU2V8HmuK7GSg5Tln9bTNPHiTxsbUaf
iKZ1T6ZnvPHgyw+uhOxIRRvnMgth8RzUqwM0LS0jdIAt8C3Ee18JjnSc64XmaFgX
zsJYHdTVNBZaU349gd9tkjdevtkI7krWM6rSDmOY8ySNlcC1+F30p6ZU5QrF8YD9
Ysj1Wse8E+n6yywCW+aRhgp2AJte2rA1pkvu3EVgBX7S0P0HmxJVoNf6+jeCwCC9
R/e1eLedczZHte6raXvF3HRBY/sqHLI4aanXTCE8zNB8o4d3iNi3dRXT/Y0Oqnp0
oOMWnEzEdD93MXzUTsC7795RQlj5vT6sqGGzLNs8921a9Gq6r6kmNkDLmV00j1S8
H1W0hSClFVgglMCJL2M7oS/vgSRImwYWZKIMjxGiStL4nUw2t/1Cq81HJ5X8EZxm
HMP5IYtM6R3TcQm4b1fcQc4iWOoQsp4Flz1yPpbLO0DVgA6dByzOayAZFfQb9YiB
PK06WzVofrEAKlYyJKBF/Pt7uGCJ3S9Oht5xE67d+xrC9dqhWfl7IkQsmLrNx7ED
6e/tPXTv7gVH/AVgFq1BTjuVEQtZ/Q0saSTev1Tyi0N1vezkgjCykTlG+T9tW7hB
4H40H52I+kNlUbvMakVRcVMvQ6/KBnwR0cWsEZFZcGmDq5E04TkHKebI3nwoVv+c
wMdVf2P/uPhMjYzgKYo9Cpwm/llrXAfjreQGdl1oGwQ3Fg+tQeNlgso5DywyC7aW
yPmETmfFrz4fpbEPGCcrJ703MvA+jXPPn4gWqDMU5+c/wR3TWZROG6Xz5hkE/a45
mCG3pBWlQbDpvNwxsg7Q2SyqvHd0frFyQnsZ30e3sda7aE3mr5XqSpUSoG5IdXVw
Ii9519ko0xDf/kJDBxAGauS5jbBjyf1CNqK8i1I9Z1qGHIrPk9/XzQFS3wKsj+pA
QEoyg+vfHjbxKp6pC9NfxvEn/pESV5OVWP5nZKVidRzc4GMeFGG3ymbBBm2e7Iyx
VVgqAvESC6YF6TnJtHZR42CYT1fpedo+ZwZi9im+S6u/9QQLotTKIObqOQUMCD/a
3zuonIc1Wn732pNUw6B+b+K0oiinBvuSqpW4/z9mWcZo3yv/aXjqMKKY12F82OhG
Mz90oPiiyDAD4ljeRHQSUdNYYEdt0PwljKqgPDLG4s9XRntkASdFwHQzxOWJY+/3
R7Ra5cuRYcGkzEcUckiZ36ezHab0PQ/lznpNiN11X/lAhfIO1dP71qrbTSMLisbi
rSaY2T6Hg87K5T9Xyg3Zi9BdnmSv4AiuxsknF1m2ZSbhqCnfpHHE6II+N9cbaWUW
xbIBnrLomnxHsW+DaYNnBUXB2MyQIp7DxzK8GXmED2aJda90FMeixODo41FA4eHI
aFJEH+iOy+BE1M3F0mlkBw/Yob5TfRe4rJ5daZuorbgVBRLf33w6VSgigiU/GuUo
jmB2dTSOXVVWT8X08cqLXUbzOfuyNXuJp3M9ibcqpSoPy+BP5VEieimn7Hr4WqQr
6npNcPYbcAbKfmB1qsoTUzp2b+qs2+Wu3grt23VsusjIvJFZNbkcAEg2i9sCYvPA
Hkt4QQKZ3Qhm9/H6LBs6EBAY6nGGTTub6Qkt+oMrQUZnjZ7BJPZykt0wmMtS9Go3
XnmbrvQa6ju643v2mhG40CtoFVI8vvE9cOmwMrHarGTeEFWjF6uxZDLt3gmSb5V0
PX/GDCbS9+EXWBGmsg7S04+NST27TrmJsTO7E0X8tvqRN6fOrUUCS3hqhqhlUt0I
61Yu23mlqUKGXotb2u50FOq+U/RVRPSEHQrdF7ZnuK+dsWETI7XbgvCpsFeD6ai5
OnsxzT0BOaqN7sjgd8CrTHVUSQAH0NvIn9H5b2CA7k4Tvv/HSBxZtHv8Td/dZUHS
wF2soYs3HvG1+yOYValCpqPWErrdk2OL8dY4FdodULfXleKi3HKrG925B4Ps000R
0jptYzWXUJLTwzP+m3ACZFUNYV/NsiGHqEvXquchxHNzDu5bAS6z7U8UVbwCiTIa
7VroP/X2vqHAyfKMp60tUJB0aj1H/N3P4t+GONo0weY4NK1lKqyXWPxoq8SVjECd
u2aaKENvZ8VZZaa7v+5G85gJSQ5TAFJuxpUGJGxyX2Wq7tZdinVRzP7XynxbP72z
wsFYckCFCKP9a5H6Jj3Z+JrdRLP7IqA3PIPfgbBAih9ntg8MnD8GLVG8DpRTyWPc
WvsIJsKjQUdnM8Z6a2h8+RWR59btTfDcEtMEhUMcla91KAUZJR6zMsGF/t6QySqA
qEM2LsMaDdT4m3rGmmvhVLXbgmRULtuLFiX/0pgb2XZMXDlXw50Tl7X9LJy6wDr/
91m30O4gB2ihqGQ/8GsDdAcuIK/8VJwU9tmGueNWCfsU6pn47VxOxcx1GGYfL5HG
0ABOflT3Iul3HPW2jKuwJg3TEIZUF2i34rwWMNA2ZqBs2baUc3s1iNCZ3I4zxFjS
fMvgpiUYlI+oMN9appiWg2heRSVU4+iwfqCUGAjH1vJKlwlEgKrDHTNlYVsq0Ns/
bQmnBYAUNrRoGVZkw7SoTIm2RYRms9kfYLZWVxZ5IrJPDN0NB543UYziZrU0ObAv
g3SiAtgF/nIyoHw6LAIyo1/NVpolk53vf8Y6wu7HIDwC6SUd2oCExtAX73dUHdvC
H+DQmK6tG1guZXKuZ8JcB1+qGfb/iAF02YEvZhCcb1yNqehLz6YFLtUER6RkRnXF
J2Yo5+9C+JYTsF08uiP/u6RqaTtSnEsTcR50VHAMP/uuyPzLFDscirbWmGEE4wFx
1D0WAGghZuuyC1V7Ugg4phSRmW3431RJiRKPNRBmkFNYguFoVDKvWqmlX60eGWQE
l2QQw6olxccxI/6aNW6vQ4q0JV4TpPBr81jXkPf+JTb9oWOTbAI/6tPlHC0Ewrkp
xAaJpn9CHuAPQ52B0uePe88u2hCbAwGC496tObFtuPBiLzP+hT9Ag5IhTI48/cmf
0ISnWBi3B78tt2BELetr0WQ6SK1vxUovEA0jt5jgjIum35U5kVdiEEb87SNz9W52
wq1H44+gGzgDBm8G2fhvJcuz52GzU/inO82a3pzGw3t9Sq4Aq8flHq10e4A0Io9U
HdCcN6xQdtPogECzfobeRyYkuTdqLYutJwa8ucw52kPQwrfabD54l7RAyMqRGrHD
tVBrBWpnNTrS+yJta9gs876zk2CJuX8TApIZ5ihIIuY4RCyeAPp57E8AWdF0rOKZ
gp6kgLm3kItZB/zzjFZCWDhzQ9Ilvv8LS0KeqqRZP/Bp/s23BfxIOPK/lByhwKd/
SKHAugNimvlygS/YaBkJbFFxA1yHKYI4Y15NdqiAHw+XauXg/sJL9YzIPRQCdRSi
dycNALwgxBOVokAtJHVqvWHtp3GekKJGI0n58s5a0SOGn3vnxaYVeMFtzB7m2sS0
fZYoFm7bi18E0JuEfgEDeqEZG4vsBI4Iv2jKunxff4UoX73Osi6lANihCkPkq9To
ZXJqVd/5KlPCpqlsXn3KUD19qqBZ0YM0kb7IasuEXb0KQWea0CJvvxphUQHX9XPu
evtQ0CG9MRdZccY4iMuOIc5KOcS6X7KbH/QU3uSx8yVb2A9fryfx353UVr/5CWHQ
uZpnSWmi5HE55kb2q8P3tNkEqFx5QEOUm1e6tJaOujmJSyHNIYJm4dfTw7gsvYbN
Lex6yWCUqYZvRbQHVNUu/9m1YfLNPsreMbLUhyS0r64y2PfEvEAHsHRPELXPp6qt
vPIZChNdhlthfMQaS8ok2GG2fY9yvCgjw8TpttBsEimuFzIC7uY6nmw/SJFGzGcr
nSNiprwzlG8ZW9tDEz8ldg1t1b0I4OuJqm/JUE15QrPxQS+L7r7R6fIm9hiJeaVC
Znk+boZlBKHe1t3sAtuneJsoijV+zQn1Rz0W7Gi8ttqosL03jTNsdihdLERd/3OC
/Tby5y0aRJmD9bQBfxXRWvquu+avijYYLiULWATHujK3X46t3etFL7HaNwnXvjcF
ui1T0wk1vNDy4Q9AnsjvECcELCGIMel+yFOVBXd8nYCj0mZI+bu5O1Lf8r8LY89j
D+2gP7umLjqXH5oMvC+7fOd5EJowNi3iff0MW48sjzgQRt1fX1JklpJgKWGu2GV5
qz+4C2vrzEu/XawgfPZOkJugTgXOMuYYS6GIaG3B0+IjSriMEj0i5L+5QkmhGcum
022fOQuB85a7cLq4GopAO2yHZ3tDnp+yRsjfQ0vYN0Sg6xz3ti8EIQ1uEbDLCjuU
n2E9lZRKF/SONVSeAR7MpazZObb0IpwIHkJL+N18d6ylQ1h3ry6IYnlTi7Ose1sL
UkIiT0dLG3IIsEQwTG8cWbFuoOm36TgRhURbkLmQND4sKzakz6dVXezamLR63qvn
JtppgB3gzCl0r6suVHk9+2Km/UGNd7KEaC+NklV9gQU7t9PWGtc0xHNUkOywljWY
DIzhma7f5bgS5YjhEVP0mPM+Nep/5WGQPZHaawQC1v8jYoPA2Kmq8Qtcg+ri5fPa
IPKdunnEK+fpawK3F2M7G4Z6jbhbL7dJrA2MUs7OKjd/kn/P3ESRJduDtvbW3rij
xInNwN/n7D03mo/WDnjRndlcZwslf4U+CsjiPW72h9jIyy1qLitgh4tiReJlAtXb
jip1oqBMcYOmT4twKbEGM3NkMrMKFhIMtZX05BC6K9LuuyqihVTiXd1fbJAK71RR
N7KkglutizDwxuwT98q5DSILd5Eh+o0nWfXWE1rXUQmMl8RwpIZu1MGDTj8tB9ST
0yWhS7ySl29607WzwW08djxvJ6CrksnKO7kvuX+bNT3TgRixQyMaYFNyEndmA3en
rIWWmrTrPCbHaz48DUojPOq8P7DrjQk91KUZfGaiNQ4NTTwM00HoCcWCdaLGCNs0
zEoeN1JFGDMSjYj5d34juCZ+I6otfYe8FioBK/6yxFlNwXsioFaObLefJSPg1kFQ
vgrPeIgBHFnl+PKA0JkZuzBqvTYATZSGPQFhbOryLGIZgY326gY18+S2ZOj+DoCq
79+IoOtanEOj8PLIr1KgJaZ5oTmxdzsxNreP1yLQrPffQQ3jfKAsN3+pWuP4zqnh
wjJq8Edpv0KtT3SpnSbOwTdboigE0mwRM/IEuxZ/+4nm15/K28lX72MsdHvn8L6R
62UCVNW6btWeIJQwTWBSDqBY1WKo3wzLMSBLMIX5Lc5drblyWLPXfXy/fDlnRQa+
x2LTGDRoXU3hoNIjTZiTOYw86Ctci6GSGwefCxtB6xXUL7u5Qm/h7Jw+MNoMdKdd
tQkQa6KB5QO6Mr0Km02MwJpeE56jSqRP5K6DAxghF31HxcmZ3pDpVDptuYMBG89Q
6n6h+JI4VTl7FUIzuT1NR5Bycm3t2y7tcWSK9FIErwdXU4JvvLlJVVhfuZ9GB2Mh
6q/kMMLCdgWEJ6Zv1EoLBd0SZ9UzyWZGl/uEAhDf3kUBURHEOivZUU8NfoKBznRd
oOLdE7eJjJAmUKFUjOabhHcPPnXz5YMc92SNP4qFWAUUK9DlmvOAFRO9EaS3SYKS
i9ErFp3c4njwd1cs31zTsdFOMUlegGBWEwUQRvvq9zmOqpR/Qw4Ou0smokvskHV0
F/APqzAx4zMHVh+ZKd0HJAKCMv6+2jV6kvgYr1DC1kMERUsIcr5mtYWSrflDFDAT
7GOTGdXoVBuFtKM7Vb2ZF/UbIrJeGEqUMfAzfsNQIbSyTsjE3osUHhzYPwy4hUHg
4HD5jrZqQnBPges3EGOGBr1NSij+Bo1xnmcheRF7dOqsqVkGxFD4GnQFfTAQhQOR
P1CwjNSqHKqgoq+VUaAIChBkxLnWxxGfHOqgkJSGfuAlPeFPoZ5uW6YwXbvwnJPz
Vx/N/CLiaujK+lm/aAmPbAlrHILnoVGaEFgZf9V7DQOPyAK7gQZhDn7SB0o2ZqRy
A6U1kZlWaa9QoiSe3r9PH0U6G25F8m8FS2vZuoysFsqNrDgFQFsVcEGw3MtXmNSS
fp/K82eQNkTQG7Z7fAnqk1XiwFnhRMZV5oS2k3z7GM+qle9GW4KRrNFa9mAS9aDF
NyyXmEX+8fMAKOiIsJhELObWnNcG7Sm3qp+khF6XYBTQdGQPrU6Ac9GOQUU8Catk
T/OSLiTWp6yEnmsAuGdWZwHAo9D78ErE+VuF44NRCmD8MDQKP9u2F/Ru80myOo5W
vvUxvQTmWOBa7BfbO5paUj4r3vN0L0dyV79Np1EcJAsQZaHcNw5V46Jr0HzCR1Jx
YeQTYQsMkjt4eeUGt3an6pXeVsU64C1mUCuWxryArnX6HWkGFLeDbsI669IoPBCE
skrxv1a40AP5Qj1iguQ5ZMafbBoZhQE+Hnn18Dfw4QDC8aZrVP1drbgsqI8Ux98S
KH2eqm5t2tFt8TI68pigvEyO+FGX6ekk117rWXEfsU3d/DdH3z6Mu7boBS02x8TZ
91LaehVZZsiekSjSNwow90Amu1CnCODSYz0Hai88VqLQ1J9qsj3QXONLLXjiK824
eKzy5NAT33CHxSl8XUiD3du86sK8SEg7lJ5kGuyj5GblC2hlx8HHgiP/9YCuBxDa
oqgLS6hgISDGtcjaxn8eGJ2XEnvxZyvQ3ls+UpLo3BiNeaATHQzNLN52EvGN9BBX
43cTksVcUGzJRdg9o1XzbFHe7pWt3Gouj3/NI9UhxkqNbhRuR+JYk3wzycn1lSpk
aojFzwxBneS1Kmean+Wuo+JxNR4iQg6hB+YdSP7kjlV6Y07YEDspXBvR8kHAFYEY
xqwSBMveVeBbeN2w856OVme9QqVKgYWBWngA8KLdtde7F5++vWQMksY30/sB3gp4
QJ/HjZx0jV7Yx4LEt+ESvoKZNoXIS+TIguZjJorNdIwIfAfM/bRdc7hzwSC+LfsX
Kbo9kfD24tBg4Fje2ZU5oi+64Zzc81vATSVCbKytJkyHl5+/uAzlUbjL+zGxQEIK
0dbxHkczVzDvXLHBdT85+w==
`protect end_protected