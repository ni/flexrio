`protect begin_protected
`protect version = 2
`protect encrypt_agent = "NI LabVIEW FPGA" , encrypt_agent_info = "2.0"
`protect begin_commonblock
`protect license_proxyname = "NI_LV_proxy"
`protect license_attributes = "USER,MAC,PROXYINFO=2.0"
`protect license_keyowner = "NI_LV"
`protect license_keyname = "NI_LV_2.0"
`protect license_symmetric_key_method = "aes128-cbc"
`protect license_public_key_method = "rsa"
`protect license_public_key
MIIBIjANBgkqhkiG9w0BAQEFAAOCAQ8AMIIBCgKCAQEAxngMPQrDv/s/Rz/ED4Ri
j3tGzeObw/Topab4sl+WDRl/up6SWpAfcgdqb2jvLontfkiQS2xnGoq/Ye0JJEp2
h0NYydCB5GtcEBEe+2n5YJxgiHJ5fGaPguuM6pMX2GcBfKpp3dg8hA/KVTGwvX6a
L4ThrFgEyCSRe2zVd4DpayOre1LZlFVO8X207BNIJD29reTGSFzj5fbVsHSyRpPl
kmOpFQiXMjqOtYFAwI9LyVEJpfx2B6GxwA+5zrGC/ZptmaTTj1a3Z815q1GUZu1A
dpBK2uY9B4wXer6M8yKeqGX0uxDAOW1zh7tvzBysCJoWkZD39OJJWaoaddvhq6HU
MwIDAQAB
`protect end_commonblock
`protect begin_toolblock
`protect key_keyowner = "Xilinx" , key_keyname = "xilinxt_2021_01"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
KA9cVevs/0fyPmeNmim17AMCVKqU9BLi3XLi6sBkPfg2MPuQ3yH/0ZuxdfA470z/
u54/MbaohlfCNjUztKX8uh/OshV2P1mr6kLbI2U3DzVxxNE3QvB0/bOLReH5tfCA
HwSp0e6TCR85kkGI/HgR4cXz0EbYhkdexeDWFBBJftUcmK1VNoQiZxre1wIX8nBP
m0e+Ki7I4ALlNyXGt/hU2PrY4OmWC5wImZB1jih5QRQKkS8dXMsi858KKhUGSqxY
sQxVp5T4KwqY4fvqcGFb4v9IPTv1PaKKL26MFtrgzyWo2COGjTzyA9BIrTUTUtuO
XeJqFMW4hX9VeupV+aRp7g==
`protect control xilinx_schematic_visibility = "true"
`protect rights_digest_method = "sha256"
`protect end_toolblock="B3YNvCssl4wtuyxkxEE/WbGSszv22Nu5/Dk6+ZOULiw="
`protect begin_toolblock
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 128 )
`protect key_block
k4ag3TYMGgrSuvellzxiL0xVLm7fSExLGPrQiVAIJQjOhMB7efNsO1toyprwMFky
lpUdO2SFDcPPBtqHJnMt1l4pzqeGpxb9ujsag+NS3MY9YgQjc3FBgfnhDF83xz3F
lN6qXDpBcn3SMrfJ1DFAaxEZtrhiJ+oCBmGuxnjq9C0=
`protect rights_digest_method = "sha256"
`protect end_toolblock="0ekDx/VTf7Cegpk27kILstUnKeU0jJYj82NrNmdF4Vk="
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64", line_length = 64 , bytes = 16560 )
`protect data_block
u06ItCWb1FF+sqwNrSG9xyGjK7OjnGLyDHAWX4ImnyqsYLGqBN4FCzmrHPkcA1tf
+Z3pWW1O3Oo3NTarqZfZ7zGdNhLGQ8DKRajAeBHh/eh/dq9R/IgVcu6S9fhL+pby
S993bpJjwxtMDn0RNN54X1MSvtEYYT/sbwehd3VbjB87d2xXabFNseJguD0a8E6x
it7CwxbrNVcl8rdyQVaDF+KjSglu2UXKqRcZ0vMSHXy1ORCbtmvCg38SlrUeLF7z
eoc0AQWyqowP7RbgNAsn55nr2iqTK9uoRrOXOyeN/mVhwThOzYwwmuphE6Ou+6LT
f/QqdwqXQHDbj2/z2wblB6nvRG/HZ7YLhHTInkwd+Qlhh3ysSlVV10zLHLW3QMqH
bwqYtB90mTXx/YNXRkTXAisslReXub5xo1aCCrol5y+3n+t3ChZVCs/q3mD4gndN
c20xk5OWHx+GLEsdoBrKZdWOIhmiwkXeKa5IvluV6A2RObVNmDsL5+q7VmkiM6Pr
Zbk54uxZV7VbeHISKnPbgq/9ZeRksqXcgAyhQE/A7EhxAHcIITujx73XBEpvasVY
L8H4+6PFCBZOpScO68qLbDeUGPMgDKRtgggTbaUQ6qlVDsXC0mj5GeuinXz5fxfh
c66dOn5wVwJlbnWfiOg2WVfk71bmqggEh3Z+AFA+4wnaD8ZSo6R1KK/CYRSOcHY3
ApHiwSIGdrObDcoNYbvZd6Q4WS6OcVN/t6nOnfOkSDNiQBvPbVbg94Tdv2iLNgx9
NjU5tNUMyhULSS4djDWIOo2b41iZNawNTn0eSMFRGg7RtVNS0RlIz2dmQ1Xf8gfM
94uBAjoQVvZ2C2AS52wPQ539dCcDqGHHWp2PhWPYrGLIY+9DX4fFTWyetFYMs9/G
gW3bhl1qKaciiXTYhXqzvd4WWlEmnj8iKiG3ZhPm7dSZFCQvWzKt3HbeKMoitXEl
A8PRu29YLM2PneeFa3dljS8VR+e5rOdtbm+rJAxTurTkfSK/cGhV0gRs7bNMHjFh
Pa144gLGFmN4VxRVzFjhQjKdIl1BHErBKwL5R37WCmAAOmsfNAue0v5dcyQ6JXAu
5ix2xrhB3+UDrTEKbPeJHFnzZtdjHkaYUSI7MRKTxIj1BUihlgMoQXmSYu9ncGX4
zP7RUzgrsbjJ6X/GrFoMlslegz1Y8WZRRMmAPEKc449Sbp2zTCgmiBVbRSRBrpYx
JQboDQgZ1guRzn/NQGWdgBYUgP8CPV2lyXDA8LvbD3eBitXk3snTHSbWmYqyIRiB
z/zDqmk+udnabkYBnTX+u1XiOcRtAqnJzrsvXHtaT0zTm4562UBU4/KoHMnYWAcl
AZ2Uw7SPwJUmu1U/SmjGXtlEZe0KU0s1riZ/ZtZ3qd7flE8O+4vP+A+ZHsZw2eF8
OLxZAWHd+l0S3AGmb+c1wIJGaUKVFMOPOrDZvx5jtMfqgVbZB7x87x1IB9tAtNc3
i3p9tZXRuoU2j+NM77YZOCW5ExL353NfHZLny5XB0A44CAT77Q7g0wChu/8uowHc
X5MfWIMHhgUOnwtBNIQXzTd6pxgCY+yYtbtLmOxWGHseHpq61vffopDQlyLn83JN
t0TxZH7jq+WNrsqUWc25t14A5TO7G+4YOIL1cvxB0UyAoG3+Xn4V2cQCwj3Rxguk
yFH0imDJWMxyQh9V07yG8VE7qHsLf1BKkKrWObeJqEwna4xWxVaoElH/3gW47Vom
TZJI6uy1dsjaiGO/RWZLZIVZ7w+PHFe2zCa/RReASylPfM+1Sxl10fIqZn2Brs77
Zg+cIdN7UA0n0r7RGg/+qLDV9t3l++qOW8zySj8O9V/RLrPl0sOOXZJF0whntT8P
2t+wW/D2W534Pxe06+PxjdpWs4UHe/fIhLlzDDYrJFbWSr/sHqlvaop7/Lzs862h
pgFKa9BeESZjA7iFQ5wy1nz2ToZQ5Why7pZ57J5XiMRhQTeZq8UQC0utEiWsH8VS
dBBglgNHS8zJTxdJDczLuT+37eLTkTInrHV3g4EjFUbIt/51AzLHRjjEfDIfngpf
KfWuSBrjgxeyQxbKQTpWPkuuay4Rjur2NGxg5TqwPmSJRI17GRq+9kdLUwwR5bYe
mIwhbE+Cn9N79A8Jbp9goyf30oSZRWoeGYBbCE1kuiDapKCF3LGIpKXBBV3cQMwT
6NLPoa9hYrY6f4ahp38YDHBsLLFK6wLZh7UDajKtVM1kCU5eK7yHB03W0BeIkfmq
oNGE2H500gOarBNLs/YR+ghd04Spk2WRcYXnG8f899d7Ww5algrDKVutlnOLd0Y+
hh4sfhMqIx6Ep8iL7g7nBsGzP0LFLB9iuIiPKCsOsQ6KM9YzO0za3KntUMlo0Z+S
NEGdHzcTFG+BcJIr0UidQLeCe/1q8lxOSa49jrQX0L8SXbBY1BxICV3RljhvcYJd
yRlkJvSh3vff4zgb10V3XqYn9JByY4gTDAhpBQjqQiIBVqK7+jA7xSdJdHDIP0Q2
3J+a8xd4SqEzWGI2iPsxwg1e9BdMZqo/OfutJwDaNyLKrb0Cjvt7BJ+f88W2zydj
tZq+03hd0z8BlsG/MH8wvovJmPUEgkwm/HRgE/fa2M2zhJjGrnGP1JINyB+t2oAw
aXOB1C6EPACFhErSZ1KzGwSGXR9QaHR523FJqcDs6EplyoT6vvE0o/f53NU3B2zc
VRKSS/f9xYZUcJ1oR4Uh8QUdw1dvzMDCBfzBWyGmQooBRmyaKfFsQla2pUV4CJy2
wFf/Cb4PAkZjHM2G97wMgg+/2vD5jtmknRuL75nzp5jrBTIVTnV5ZhUhKEat0SuU
APtjFUDofNrH7pOwlRxLP8r3R3yK5g/nkFLMKV73igN225ZS98piNm2Lle8wWEWT
PWrGTCfhyxJTOOpubUz7ECxz3T3c2xT0KlIqj4jsNCkMUvBwZYg9nFqCX+ADdL9Q
n7xH1R2fn3OLpRBGowearDY7G8/16yos5iM56rBbj7nmae15krolAGH5acBkS0b2
q14HG0OuoHOhmdBkNl2IdIl9d2Q16RIrlvhcgYH2nIPAlxMULdjDPuf3NI5DUsae
XFfOBR7X8k8/b8Ps+6h6iLNg32eedOLSVnpB3/SBO5L6SRsAvWp+aOiaXuZznAHH
SmgH4sDJJu09Qkjvk5LSTQMCCkChAuOhtgjGbY11yPcvCtJ7bvrOsH9jkjA7gY1C
WqUHUNc9qs28M1IYtQYYSy1gbIGnvuOiBUmJmTVr5K8Wv8B8JRYxKoCth71Gwbze
IebLhuhBD3pQj+ZUV+IyTiUCLgR64L/NRl+jZ29YBj/IsGnf7bD+kZCmo5R2aIf0
bqXhuWLAOBW9gcg9vv+17KrKskHCQIFtZV9Z3wvRKVFW/mcYV5vYrcvA5XxuF5PT
VYTQ/wRBbzFjyJJC36Eu3Ddhae8qBEzRWYerXIK7zKQFtyJhHmYkty4v56IQb47S
K4LQN8lld/QMFakwj6VzTlS+dNiZz2wpezopzfTD62hIv4/1gDzMGGnCxLLIT99f
8hFviDkSQYW4Yw6rQa8dKBT6OrPnih6yDazzMHi+gPEorwrxTUxE47MGfoHBAVxZ
sHEBXYK/0ox2BX6XRx+NUwVhRiZGjElcBWXJHtK/ew9maifORHucf6th80KVh8wJ
ciWyf3s/bT2yQ0C6FJXTtZ4mvaIpTOtO0Z46qmFFyi2PEM3D51EYqZKfp6I2BpQj
MQ/KKP7zCU7H34IS1ptSq/4W6OpEB+U8IyzotJYZZV9IG+2VOMX8Og09A7n96JQq
vdP1/m0D75nCHldfMiryBfgnm2py71UxF51YSF0QOTf3aFXl92oK/xqlWnMIAoNV
6RKAc5VFkYXLWfpqVRaIQYIQQIAv0VM3tUv/i+XZvuCzANBIPY2eLOsSX/XKOU7L
FJesaQv+PZ9zJ5/Kb7Pb/Jnyi8eWDM079YNWr7epKJtQlRyDTBXJrkz+aSf1oBpb
HAboe7ZmuWltY2irnsDAhIht48EB1iFaNfx86uaCVbSWoedsRwjmKqSqvbD6JO3w
/ZXf+rzJSFNxxllLHuq0z9jb4KRHoc1WPQC+Q7ENu5CplLtNLtO9LHOMcZDWgjH1
bi6NPvDk60zVgmWJ7i+0T1eTlGT7vKSEssF7wUF05t2p7pNFa+eJJVdzNUUXfwFs
FOJJeKAvAgQf0ayeT0Da2NaGXAY676coypm579GmBk0y5tx4w/J+YWhA3rd5v+U0
qjzr+8ccSnLrbE0By7hbBsAPKEvGDw8AwCDga624z5pWNZLZ9IS8K5xhCl58COtd
mq2aK0yFxuZrqlSRyQ9j0ki3VFi/6jMGjuCDDkqHTfbrBhvuxWeg7fb3/iN7V+QC
7RoWcIBMV2kIQ7ORtpiaddfCP02Qk3i0/H5Ms0bdbtwD1Ki/yNuRhasAHlNN5eyg
oO5npU9v3QKhjcs5MQgNXn8GYHTyOTgtNcjY6rt5omkSbqY8y7wbIpoXZZ2PxD5L
MlNuIeUdwvAnjehtO9Wjt85FaYKsRwiUXPwhKMjjL2jGXF5rP8dX+6moAb2Ve3XT
PXOWeOuzSnuUG9SjkItKh6rlBa4DaNtVUfT5UpAYBPNzEY9ePhQNbg7JcjdLJ9NQ
uZlgcKVnz3JQ1xBqf+qsjqlXxZ3+aN0eZSetN8PEOr5SwtXB4t+BiWjvqHFjxKh0
Bo7DA1/wPkqImaq6u6sji/8av3Qe+OfgPdVKfO+7YWVUeUOkHzZ6PqK0ykjdUsI8
0TVWulAQUxlpv6BGLlHe9Ip4w5BUDSStQAosfnhj7focuTFNC2X7+FUfg1UEEPOm
b+8Fe0mRLbffeK5UQOrFCiLfVUDA9QehkmYgOrR4fyCJ9vW+6FUJWCns+kge5a//
1s08ZY8kFBA4Zpzu/568wJ6g3JH2RTv3U/ontE7MbnSy+k/zbEXm9tJDiFflNFOk
OEJ7ELfGRrTn7sYtIBY2zTgyV94ccJf5iE/Zbzdz4ylWuqn7CnZYim5BnKRs5D1i
RkvY3zd1cHnau9ywKMJOWWTs9yzxDRQnJRRNy/mzHJ10n20nkeWpXT0MY+skhoJY
buAtsU9+/4OiMKNH7lDlbuPKNU3cFUw93CZB+Ve5/2oHgET/sIg3NYnhDTQVebCK
kJjtpSi6LQlYEuCpBPYMGpNCYcXVDfKzQgSk/mwOcNt6D7pMqxBMVbbcr12Wwvhl
Osd+/oovyJkzUYP1RMy9pcc0gyJiJYL8s5TgeTGCVlVzz0ESC/8yiuirT7klLPJd
pZ+il5p7CxsqqCslGTaQe5JhgTGg4/ZlUidgecWko8hYRDGjL4X/Ex1vuCnsvhtp
5wtXLdOBcN0mEZgh/+TRhvTbhVCGWxHDAtxZGK9GhSH1XkSQkt4hAKnfMJ2XaifF
VsT84rdBQpdh+Zpi2ITxtd+t32b6HOn63jGECUfz/bNeKZEcIR9XcJdAUfLuB6ux
pJtQj7zCXB2vjsF1CrbUf2QDpBvMIbiLUDfSDnSRgRy9Oc5E4CPD81/ltFlV5+yx
paWGilbVCXUeVIbpPuYhtdNZQBT3lYhgIx19hPAwplVVecBn20eGcgS1CHC6ZuO2
uT6AjJYcrp3xPIF+OxVPWp5lgck1u0MTz72y+YTuMXWgJHv8qjT2q1yMP/4wbqxg
sXuDa7ifpURBVJRbfHNbVTseZnLS4sabNkZ28YQIu11bEQ8bTCAsxrjXlNetREjr
soXqMp25VS+mG6AuHtz6A1dmrC0K98TYIets/czZOWntEJZyA/qQ44xs1hXTst82
g4y9OJ7f4fZlnkBFAuV8YW6E+0OSUYc02S8riuB+XVknvOFGFHyrbCkGCVbagW9X
3KfGcdkftZqQaYy1JQgoyByAHPIpb1vPAhPHKCk5WlI3+5S77TEHx6MLpuqxLTAy
SwGBkC6tFs7rxXS/hXO5+HFjz7wcEpB5Z/TqCmeD4ocwO8nJ3/CfpEcY33ZUIEDI
+h6rt6GwSVFYKi3IzQNUrr1FjRM/aTV7dyo7TVisbR2ZQkzl0pWej5IoXTIDU6w9
QdxraQgWgloxbeLidbwkUcgz2YjdnO6E1Zk+JuDP1KnvoPflYGGPd39MO0bWIQWv
pW7dg1XliilYwYmgNADa6uCrNi+4x21BcsnIfZbxwbOANROi1zxNmtIy6rXFcV6y
g32nuXtAHyA1L0t79aYs5bM3Hr9VyLlm+2wwYd9Jb5ZcgEgLjG3etGXkWLUSW6Go
Wf/R5bNjKuhafgze+meuqxtXvr6UTXRuxLFSQ9v11ZaXzHfwxotuYYFv1BdQQ2j0
Olj9VNYX3h+SwLQKTBm6jWElhcVJvm5N7qFrLX6/gGsypf2+Vwi0N+RHuVQrjaLO
Xh7P9njBRS6nG5hX2uM3ZmVAG03W+duyy99r7DceK/j6EJWShtCamtvHalUJEuDO
cZ/eck0MvbuVWa9euDWjYErWFbg0cg8oyCj5WGaQEQkj+BsUSsVbWUjPYLJE3AZh
bVBrH6yVhjE0JSKwgguYAye3aHDFub43Ohz6cHSGssfhZl/oQkeiQZY7qA00Jiij
PFB5keaSNLxhKuGs/+FDDKYL//DFgTZfG1xmEQQ0O63AREoydDsTKf67Ud7Zw1gK
iVQ8EiBDdX5doxjKpqGSPDixU9UffGr4fYrjVckkAhjDyQg+COWWmmD6ON7YnilE
Kjuf7sBZBFrq5apVse5Q/RfP9YPgu21tcCXZCPHSsU84ggKmIT2/45P48UlML77w
hC1VDB2gW2V3gbJwjE7D1bkli9anaqucKSXfb1z4dBdW0quePC6qqvIZnUkYglBk
ldNcN5f9L4v9eMEMeAKkE/LQZT4N8zGlDJu6UJT81oxKlIxCDF43uUgLV6HhOzhs
kTQpchsg2YzH23288zPacg8N8/Ixcv4zAnyPn+Xl8kYIUFJNJu54sC5LxJb9sNQB
6PnLtMCeFd3hKYU4cpbh+u9lI04R6ZvTGg/351ipVEZnfgqmO1wnlGhBnq8VbMIg
sngsmXv9tNpZyLX3SQOXzpIrzCDlyR5RYsC8xAYv6xIU0CMxPVE6S2xkmTKlGnzF
SFzKF9xN+KaVKR+ykE0t+PLj92XjkVXBC4+VceACOfySze1GZWq5rT+KyeeA/LBf
K0OvOQaxUdx4ibQn+xgr9B84hNJk17h6b49ZIo/DBhWbNCo3q3wSPSGcpypMZmNL
2rCqYRrDmz7hZhh50ssN2EJ5ih0eLpozKSr8bBWGUTAbV9QsPJ7VLBwBQX8Tn8TO
WZvuii0z4mpTAS/5SoAZDWOlW1GysP2UO2VJMLuK6W8UAa5GbzW4v+89cihAMise
PdITdA9XUN3kjGlicvKUQawlzm9IhY4Z17MzK+T9V1+kYUZkjstVSXE57R6PcQ89
rO5bwuVkO0x+qZ/BIaUMhxm6LaNo8VK8UgtVYk0YyHJinsZVDPvhyxMzaXndMJSS
qnBSwMgnFhriFnizhEo1N8jkTNbyUWqQs3q4GW7W0lD/f2e+4q8qlzOPcSSYGFm2
HSmrzkerf5dWFmdAp3C1TGVZoBat50DbXev8ZH3smVIVpNrs2YWK74FRT05KXNSh
v6bWEL0JCPwtpdqbKNQGUkNJaUOgKgvSraImiE6Mm+lOCramNfkRmBxTdAGM8XCV
FMcegBT+F49O5vyjxfXZnn/4AAr4oGLvzMzTYUQzIq1xlO/kh0l4K5+9oHvgHH6L
3mvWndoxV907luu08uF4WbikRSZ7usIF+HmVgBOFTONF+9B1UwS7N3hNHF/fBD3z
ugTTB870P4QP3z/tTV/GWIXt2dtRL3YU1t9hW3GI+qHzrOFeL3aQvkoWHLpO1Dl8
HfN60eEs4ZeDXlUu25A5zYn7xJpzm2ZucIrTU9OFC5RXf1SH589lETZ4r7DswhC5
R6mi/L3Q+z3pDv4K8G8UF/v2mtcZ8Szwbp6H7J4EmEflPDR/4Ngtxqd8IoODJ4f5
AS9WhCR4PyTR91cUOSf2CzDIe5pp4Y2+C4IV4HvwesDJiHEoPwbmQzl/RN5pktXr
d1SRDi5X0vCC5NDTGnSVjFRbsoWJ8MZFt1AzDtRckI+fEEm/kj3hX3eDoMJUxqJk
BBhIVzyoFk/GNiJVkSswCX62y9nRGuC5zPDRknjyk9TzD6pn0qcek0IGF1t3+ipp
V/2IgP+WDdS0Mbe8vo89vwdCmmeEK0DAl0b/AQm7IYeYjuZxbpGEBBD8j9fnUtAp
dGe3doHIARvlntg8M7Rc1UzJrcV4Am3n6Qps7nCXevkKDBxHqDHpr2tU5WZ+vHoz
s/7vuHK6vhGB/FWxsG9rGi+tWd1DrMA+1/7SNB5xdU/Xu9CP6+lny5HfSHTLBF8B
oZDtD4wzcmz2HKYZ5U4HTCBJt0fCKqOezRJNXMNYLCcqsiSS4LnrwLP4YwieXnNN
2cOJS4+oyOa0nCnKbMrECT4XpODKagRnU+4wBUDJCM/SY37ITCaVMMDpKjj87cGE
psL4qBNVRGqiloQGzjicyzDqb+WUoIkj3mfN4ErUIsELq8g4XgoDFlJRZ7ilhWQR
7/ftcfPdFhH5QU9pDh8CuFUf5yNgzFziMbDJ0A3vW0YUR/ojZTTk5kVhc2N4oKpO
5tUv0qXkwSUr8rBbsyFHUYt65liLIZRWB9Wq7yge26rx+DK8s1RXLuJT59Df8Nor
7q750hmO70K3kyKANjweybKQeCC6WoGw+McQavn0fVQeyQxwsaQlM8udpEoTx8mO
drIXmEXLgXwL51a+pkTnsuKluVJ0RXAQtqjLYI4E4sn1js9psXSIfDEg9mdOmOpC
uUjoULiGQ9Nahx7mskc1dictE3BC0uQtBpvIce8KgszM+uvQZzRpgRJLTTzPsM38
N/12y/sl3tHb63X1Tid2Urx5gPxlwtZsU3M/zFbuDSApLDA4UUpGNWAgJicgqLfb
sVd7xjF3xH2Cj4t/HwdxixcLHFacBdLU9Zbwe9tQBSZ/0W0JMtafVJWqCHQluMuo
F9UUIa9+zGusUQSKMz+hqa01IFk8CgIrHNMPUSTVpu+BqZ0R+1rtcNOY+VmXoZqV
g48i4xrioUOGrJO8/adj5enB+A8zLrdr09629yjThh/vEAgK59ENzvTiiYotxYWx
LU0FCBwVPsIcZoJ0tRNn1VjrHzvwTkUMi47E3FGnOf0nYP3LdXNZcoxXgUuOrH/K
I7H6f0LuDoy6D1g7n2elySohuHiWYAPM/lBL29Asp0wTr10CY4rIq+vZAooIO7QC
4hFRMHZAv+odwabWFQ529lFZhi2ghGKmh4l3f/Wh7F8HY9R6u044RsgTkO8A0CzH
DiPhOXlAfx0aGnOsxjk6jLtgAV7njfb0IzMTdSK5s7ExmNog0pb94PkJ1GX8kNxJ
xRznS95XIsBGNagu8ESJCgI8yV1sxEBofyBMu8LitxPoUc4T7n93M7Ke/C6HPbyB
1oUGgInR0n583+e6spJQeNCJAa0uG+HOHxUEeJvAilv6LM20yaRRiGEbNUPWHl6i
hBl5jonjvCUO53REXuNdOHvZ9rKFrMPwrsDeY2rJAsy1EF6QuoWgyNqCwKg0/8kr
uQbxLEQfczMkGRX5fT3xj8B2CTHaRgIdumcJNFDx+IKDNJTq0ukvUQ0djciE34gD
Qms5OpfwXeEjk8ioxj67Gvaeb+/EDoDMGPhoKYMd2NkLYOMYRYStoUt6oTzQBMe2
rP7QaPyrWqPIbW1aIO5+Cb6gMdVVOaqmefGNrZ+NoSYBEwoKJGpvPZSmW4C+qe5K
0HabzXqxPkvbQVOHYpdW4EliS2kaufBIbEC0WXF7lRflqA34gjli5Z6Z8X8Mz4FK
p3uR7+VHHC9h1S5D76pIhciK4zvrm/63Jn32X7/6XnBdty7Ry8CrZhZM85dDwtKZ
uMdvGJR6hbDht7ISD2jt4IeI4X8qoK3pYT13ywzRuKtnzphIpfO++HT6FWoYY0Gq
TSP3Ltayfuz+Gc5chxTT2BGTF3VCAmqcwpJUAX7RYLC/I1K+V3ln8y8kCVJExFYZ
Y8mequ9sEnORLPf2oi9p+bk18sO7ytZKMiKP8v0tnGOjkbAUv6WIPRVx+obU8bFh
VIGOQ41SXsavqIvnYokBf0qO9a+hfAU5wjAUPrkB9KsRBXJHfeURaJ6OyC+Ehd6L
uh6B18hAJpGQqg6HmKR8NPQovHzsvrxo8K0O+RW6sb5cRmZ0OV7O+ZKB+B8SuMxr
EhB6OlOtjAc5CtHjYV3sZkrQIPYirdhPRNN6OPIh4sxxJbzJznZZWW6d+SLiOm2N
WK2EDSn/J3YaW/oJGXOY1ihLM9/p7LKHEVfT9GqYr0ZYLcepSVUs/cFzEVRr4E/9
XwmiUt6qQPxyH6Uxrq4cCsLYTm0jQL0Dp/7YMa7PshkKxxp+WJ/vYUzpod3BYPJB
tTKPl34g5ZPtdqR+x9Rz+HXROKTRXFMENdQc100XMVp7lRAc2a0a2KBk3vAt7gmm
dQIZ3HiGMh0Cbx1zA+LJ6w5BknTCLC1cbggQd7gIL+ReHvPBTzTrK+R8UzSpmY3u
P/B491InGqL2lWSn/KbMc619fDzilOq8HRVZsLfY5WQn2vq82NIRgn7TmHxlGXbU
MtGjlYPXZ394r3AhsdwaIsKkLjfjwuql8dNCJHoml+wj/rnbKSoNMTx72Hgxoe9h
lTyk203wANbYVuRLl2To4+SmDsHhNr1zxFS7OLAz3pFn/qpXOIzSIOLKkirELWIv
/dXGRKtswRJoLe8rxaoa1gu/vpNZoZsHNKi+XbMplL3aEdq7sO6frHsTOo8b5kDx
tkonRTeB94kpL80SK0bJ/rw0rqXw5/pFx6sMOSM6fDCV8sVANAukqiJQh2ahhjR/
/2mJcKqvS7T1HmOryo6gTJlyJszD9vu9M1J+yjUwZtJ+JBvx/dozHcxcWOynV43H
Sl0rqH6sUZUgRFU7IXOaFvFokkS7Ox10zV7bCBel8DP+nOTCkzxnJ+oiml5TPYXH
lynIZsoOyZKsBLXeaQX5+emCZUuaxOJ9JYb2ZCyDrCT+TvQs/2jmO85NOLul53sK
DRUOCRmeJjEklsmyZRYg4aGqDnTzjnMGmib75IdOXro4GGGiBE9UBTcMU3kzlB+b
mA9p53IZkPR1bv7ZA8SQak+67a5VNhiYsXfxzAlBi6uulqDr31oruerMfgpydSpD
SdVHoAOrT/wUoWREoOMtQomxmC2VKyL5T3qEjmFvPS1fqNccHKCJ7lKUsWcoQXaY
0O+V9uUIzwZcWtX39EMN1hsnhD2MJGRv8fL/hNH+1FlusH5xiqUXWQzraJ4kpMK3
wUz19AxB/Xc+TajYbo97im4LGQfCm8e1XffMO+Imjscw6cy3R6zTICNRu+47jyCs
vSCxuBNRz8Wc2KM0P/grbQ0TiUxbK7mnjagIiyFnI86beO9vBuVw86+7eWbP5iI3
Si3BpSHOvFQBbdkoMLqQ7zitHnw7w6rVOS9vZwaxGaEbEsu5Psje0grDck5VcUbE
CdcUbr4na0VIVWv6MmbB/jWRIfocv053XrzS04d9WpfEx7FyuSIu+RL3hQ2mNxaj
2Zo6WaYkmy33iZ9idiOI5GawLrfTbsqtw9UR0dPsN9J1P9RKrj+Z0Tsp/59KU7A2
vrr20CRuGZ9XmgyK/oEfxLbyJnA1+HVT+xUgJL5dyO9LkLaSSKNusLqw32uybGUd
94z86Ii8TyXN8HTqFrMeq1w2EzTnJWKugSLfQZQYEn3GVSOEfLOMC49UqlRILRko
eVdghoW8Xu06eeFCW+tnKoXvw0CdetJ9IORZVRv/je3OKOMbsvdbCx7JZAMLTaRo
N+HZppG8b8jvwcDpDgA/V1dpNOuWEDiCNkwrr4yC6x7kABrQnMo/F3qHCxQJuKMg
pDtyFcYSxGTKa6LNUSNeZ1uuH7Ojk2I3xSIxqGTlZH17sgVL+JoZlIiLcyRg7Nol
oDx1vBmdvlktIevcqE4uLRQrm1+zSn66l+Mkk/OAzy5ePhM+hSBA5Z0FJ/as0mW1
rMU23HgHKRifu6MO/CW3qiyl6Ief5DZDcAwKn/1Oio1Q2LuvnfQy8EPOMK8YDT/6
JQUyuEKuQp6fuRP2gQTlu6OGHts9g3bxoN0SbyP8FwghtwTI4uRSbGLYNTsYYKW6
brT3IBCe5v8zSsvBZD1Riu10gzVLi7mPBbf1TS/0QqJ4XrfQWpwZL8RxDk9lP27Z
prgsHo0F//0bcfKnY5XqIKGgbmP38NA11kn6QuBiPIX1XJCmsFiTm5qFxddFSUnw
cKCOeG8IMtKvylKhZ028Gl4OmjG7B0psP3Two9+NH7JjZ5ZQrRvtUeM6fOt2M45A
6J1xWqA7CxdZasCB+yq6TDKHo6hi8LutkrT+rvTuNbBORp/IuKUREwxlTOPdyDN6
VbSPsjmhrYFqG5YFGCcUA0WCwmgjgjTdSnVV1K03LOPLj4oF792pxKuDHdw7HxuN
YhlNioKavUftQpVGqPHPJACwiVIzlQ2xG30UfcozDhLQGLGNvY2IazvNLYvhLj9v
AEn5Xti2BUsiLEdjZoAlvKPo9ug3uqgPxXS2gjlfOZOXFErKEm5UpsNlH2270Q83
j7wMkTorb59f9l++arqb4mOi5zqkJTVFq0zfu7DkpIfmX2gyh3/t1a8vj96wtQcN
OWXiExCTh1E9NebNnQVBzeKxaOVMeY0NBhSmwxe968sJECgd4e/OEQb41IENN44b
kF60HEMHUR7CipAf/JJglvHI5+X4LT0gym0CAXKZHsdYmy4ZVdygqpbHZBDvny6g
cKQf/04ZIit2DGN/WvCeRufB/FKj1cbf78gJ9sTtJokpiynUMh3slNjHeeQwJbHN
H8RMW0sASjhrwrsSIkpen25ylE+XliqJHo64ArAh3RDcr6ySDQpof8UxgKAFkf3r
i9K40c/fxq120czFngh3Kj+Tsl9cjiM/Btv8f+nRUDofX55N+3IDaYoX2NwuNCis
Xugpe3sW2zA7UmfEEqMZPIlNdnVmHE5ZIvt0A6hRHjnnC+f70HzA8djbGCrf1jHS
T4EbHEmhTGBK2hLZWGyL2/GbJWVi4kvvwjlk3uMgx5ZX46bV9bHGrSkLCoVFrXDW
csQVO3EIakfI+gJyOpfHSiZwfOs2YBwpmXPNVaEp9tMovGtlO6Evy8inVNhgz3Vo
1uC5Fxp4VVtkV9rK2AiGNl63WNfaE1pwz1p/pxT7Mdb8AmiVDX0Toi2GUfHYdDxR
sS8eV9S0BcO85tHevTFBAXfbbgHXtBXbEhPRx4/maND9fHNlQDd4zIdzdjEQS4QC
UkMGn122eAeYVP2kjhfXFgSsEtmqSOHMmufDtuhk4W2jS0g9XGxnohfCpNNPfV1N
Lxw+J/zCg6DHGb4jO07M2JSsmVa8vomu5xYTVLEjRJjnAZbbvi86pPgHsmAH0b6H
zh74igzTUPkiSKZGua86dfR2dZUwoukcgOlD0ws2DEzLIaM7hd6m9xqtYqdXaf+2
tndw0Rq18OKoMSdNRhuVTOjtyma8AC0IcXTQJKslU9icVNo0Y65dZfMU+1/heL+j
s500tR7zvfAdssQ1+o4Jyb0YApuAIyiHR6IjTUKoYOlnO7RJQ1lFGd9Y9J1XdlYG
mBZN6OQO9zBmKykHY5Xy4qUbn2argu5OQfXqdUPITA4TefOT4bCbEXTyHaRiqlzA
Kf5GfN4NOWxKqRfbkDWC00GVbYEuglGg/tSBEh8lrZKWkgC+rVo7tDvhkkLZHPy0
nyRHibp/GLsn80NsB1J2OPSHd5IBIq60RD+fXBfAQ5NkYX8iiheU/zpPseI5Jmaj
6f0C9Ezi8qVZZVOeO1t7lKfjFNik285f/vyvMSYCJDz203qd0DaXgUdtug2WTmA8
8zJs9ubzBnGBUj2mrFIxu0qxjP/KuIAlxFy3QLt9AkGJaMyXkwHPmGF4jN6FxfZ3
8LLuJZU//kzQE5lzJIC8CPrYNN8j+vmRG6XwJXwz5YP5z85nR2My2PUUKNHVszGa
6I303Tj09iw267QT7UMHwcVQLsLdOS5XyV5SOibizJBm9sqNQeRC6lKA8+7gYmq9
9XJNj7UQNAm1bQSut0Ok7spe5RGWmu0pKtXhARy6o5sahzWqj6gksd5hYN3ymMi6
SGY8BLaWvZgpmL16+9XrLujF16TCzPC4SVR12pmGTftrNsnYjJpsrrR9y52MTwam
TGF3QTGWvoO11sEm2ajc0P1ak5WVGuqNCMHPLx8EQsxuucWBSSLHuTcwaQyB4QpQ
Yq+LquBqMD8/dASbjJkdLNACjI1BUowIV3hWsPfhkMjBewwRChgcr5DEe3/D7E8P
FTOWFK8osD3WV51uI7FN2jpnsvRQPJVqyRQYK3yHV1N5ubUL3qvVturi9EPlhcuB
OKfiC/lazRf70a8eO51KkHftlGpxYNKdNOP/UdPS6sVN/n3WFvgMGHQB2wflgowh
2RkahicvSrUta3lyzMGvcUgVXOiIVizeoqFBq+R9ADfpHiB8PWLzXKeA1ul5q8TH
eEBEUdaJyhUIS4giUipovgSiSgpaW+Ci01YhSGFAxOgwIY6Pa89XA6JxSSeFuZdM
1+MmOIvKgcvmephyAQs2mQbA5mKPXhiF66WF45DfuOVk9hFywI/lSpJcIkWO1D0Q
0U8TdWZeNIGtuifd2saz/bzUTjj+C1MblyD3ECfEkujnQo6zkF+4ZGwSxw0O8he3
jQYPIKk9KT63V4DdPtU6klh9+fROP+venXUXaC5f/HhiMGQJ7vTo0mGna2wOAYOo
3v9YXDq/0fgjfpNNtcwD82+d+Jer25h1cR3rWYapU9IAftLeO3NQJRf0SkD0UulB
Dl3E/FpJfC0ugSRI4Cfe+mCir5pyiomanZj6n6nfQHy6HcxZGdUtjd+6C+0MW2Ki
j0MbFbMYFK0O2PSCn1EEUowCMN+39eTo+8RIW9XObPRe5lgPGXB88ewcDTKZ2J2E
ye5bJK2TR42vEXTP0vS9q/ZwfgftEKI5pIdWj5OQCRBXlepNnC0+RvZAQwodoZm1
w44u6wcbEXqLRhS7MRiXD9XKfsW6iC8TothzFH0o1sBT2jlBIm4/pODAvK97qkL9
pQi6wRrfI6lnpw9u9tn+A4lsDlttePLlzwsbHfX1SD0LMLlm2ocpxQzi3XwZfV+x
LyNbEingt5MqutX4i2dMSJiB5L+LzHoxrLSXNbHqxbq0xCSc+Y9UP39dxIRCJ1tn
BeugyQ9oKzKUB4n3weZY+Jgy5xtHTvdYWlJyvCac6aDjTd0TI+/wFaKBY3MZMjQR
JRND9p5EW9jsUN2XWX9oD1p95P2tF7bhdAp9JdFLqRKyKzMkUcT6vAzSEDEiNRFq
tfU30/uc0Zp4ADfgA23eObpTi4FbAuSHT98IEo6K9i8vdoacfOxb8oypyCE3H2dV
6za0Q/7mY13VIpV4z595qlkaEJ3IF7uNkWWiPMGPtpMyi16CR9UsqzsSfVVUEhUC
gajb6adfhPlf38J6t4l1B9jQgfNK3cYHrHkaz+PxoKcaqFrasd6z8pISpGpQqVFW
a+4zQM+W1GScthZK4Y1Y1/hYpmMrBvnf8hO1CvZ/lp+zvjwU58QMkDB/Xb4rEU53
R6x+P90ntf5++jGnYulXh/0HAvMCVXw0H1ohyNgIrFJm5/upiIxVSqk75lyGSCtC
1DhgxQEHT0gfXgc47wVRIPzfMfEo/pt8NfNpALS7FHs44ouRhbTq7WJaqOVa27NF
2TNGpiH6Mqi/Dbdmqxh4OLz9prkGgjwYZZqTOH7GkLWeXKWALmkM3Ltg1j4n+zlK
DpzIBlTjlbny5Un5I0HpvZsTmUpIqeVbMStgqHw1ggqZyTFxuDFuqF4XIRxoTqBi
amLb0GvkgsGIpjv8tB8xId1+lHsqW+0s1G3EZ9W/VH3SBlQ1hKG4C9eV4J6uOu+x
8CRTFB4aooXg8EcrM6gk6yqzIaVthT5jhsvQjS+MSZj4qrLVoLu/hGjQlHAlX224
UYGFkvpdmCvX7S/9jcpXH6OsYrxU+ugXKeABp2pkjbNlkhDn5ZwwVMImxcEp9Vsl
bc4dP9tW5hzcJJsNcqO6ohaKgGFzyVc7ebYMO/QsJTZ/3SSmnitxw1TYTYcxH37m
IJz19vr+hH7u9RatnOQxU57uyu3y6722Sh/fpiy4qApSiH49MeRcNKh8tmZfcw4v
vG0ZnmlXysE5qiWD2cTRH5zIO6MlvfW0UN1SNYdAkKHuhZvYKb3y1twmFCXxfRe5
u6B2jvnW3r7zGnXysvDER3p/jqRq3bJjGsYwLzsvwNtNwlNno9k83HXqaGqJ6VBu
mOSVujTTY8WZRb15nYfLLlnCArxGsGdL3lPFrSStnkPKBJ5bH9pReYiYm08BgHEV
fdNFd59OHrGJU9pki2uMdNrsD4PltsJhgpwFiOIsPCIkzwQ+WRTaxfuVpEzbRJzj
inkIJtfKPqzNMbHcGe26Wiut2uHThdW4RH6XOGgzdoMQUFCxFC6ys60KqpITUak1
/B4Nqe3QPD9+EI7Qo616vl1AQBQr/oHUY4ybxo/fS7kzracB4Wubzv4FGd68c5mj
TQ1N7Bdb3G+I6w+q/f3D/XpzCIDtlU03aGKi2WV3PhXXfo3RSWnb1+VJf7m+XQBI
qgfDD8nHtK2VbC1Jl09KtVCzqAHxCGupp6PRe/gJ36oeVhBeinpPpZFvY3uGcHFE
nOraxOsaFNWtXRiCMG+SzGWBjcaqwD6vyLZakF7LSxeiCzdexEbJwoAA6FwEENo5
4Dxvrq/WWPAX4M/1+fy+cCLQXBYVx2zjD5NpxY1alhNjCRYGFUwZl0wI0msnKqQg
GuhtiWtT61Y8bGTEiipnAhXvhM6GjlTDp9x5C352VwHIsIWUvsLZEW7bf3QOkKB2
4Gjs+3fRzk4j86tIjXkx2E97uCBTNlKUB91ngoOaEjTWAmjqD4LJes4hLUFFDwaX
uOVmiIQ/DGX+ENzZpRWzbxvlnJ/fF5KZ81jZPnmnc/VvtHyIDB1h6Z8DLHzzstT8
pOFBTliWdg4TQHtM90saXacGFFMOJD+rMJzv89cSOzoQwutoJGNHCGUZAZDdwj1c
8SLSpg5rMBbYhwqY+sNHhyZCANj17/HM/5zHgir28KD0jUEBrqdQG60xChXjGQs6
l3lunNk+AUbthfVv1TIJWz8skk400Sf4zZgtpvXUfzaflUCt/yz0OsjUDfcrTdnR
7r5t4WVfAt7LNuTjWIdjz2GCi1gKpb5ZHpWkdBTJv8aJoWuwJs4mJzpr+sn2q94Y
8Vj9V8Qe2Z22XsHFTHpc7/oaX3DuGS2ljJjoUob83BMj+G+Q3VtXvsJASnCxW77a
DJl6lN9SIWADpYGhwaGva/s2y65AgFIv/PXrI9RRefyE/0K6BTAu3WzQNOjszxOi
s1pmHtaUhnleQg4tLFlwMV8EBAcVUt2ilfMCAKEpheBoPyQitz7QoEKombY/x49N
cQG4fyhYzmvyhXAnP7efUuufKM3M3t6n03wuAeAPrtlnatr/RhrTGh8xD8dvzbdm
sfhkS2T8/eKRnJZMO4FDVAKFHSxVEc8Rna6mqekeNxyHjaiKAuYJ6vfbEIkQcn3i
fYS5ZBSI1dKQ9ESqOqcoYb/4lBuMlCneL/mxkj5LGkGDe1E8VXeq3Q57U72VzShR
OtUoBBhoTAM4Y79fDysUBlfAQOrqLk0WdpL2ZK9M+nMaGOCv/OHCNXQXQD0MXUhP
ZYFt60XfQMI293sQDfd+FmrKRTtS08Z2lzpVTD3sovW9x5wSE5OQAWdFwFomo12D
O59YBGaprwoR3Qpig9uMQSITU3mmLOiWfKqgKCjawlPOvtnxTpZOTrrW2VSkgag7
LFU7B0WzO4T2J4E4WP+v7U9vIaPRXXy4gsMWsJ96syOIQEez9xr2/S0wwM1CCEYl
IeTZI1BySLf2Du5I+OBWylEgrlpetKWKG1uC8Vak+UrYLvTUk7aYWfjPOsYIyiP5
/owpL8aMSY3eNpXDkpa5RZ+R9dmwYseEFnEtH417KGUQUhlYkY+tyZbvsiveuHkL
bB9mUVnRtLhNgKXpLmUVTZp6bFfjNtwlZw0nXChViww5VY2LHF+QvdAWTU4u3FT5
GPpHSRrXn719IuP2W5SiQAQA/ZH3BUDYhvj3nN3n9oB9q0HZcRVEeMY1RAaPH/oD
ZPirFAlvxUC8z7dw7F7XSkEQqf6ul3PSZDsrsPUnSG6Llh0VOqvqK8S4LkDPoGtx
yfsxp7lf/o1ZltTfsj5VwQ+XYABkURTrI5YDD4CnahcjkjjiB1lvFP8ipbpZLjeH
VfMZCYgN2AebqaZoqr5Ykr24TDOrcBIddqY+8xMpCEsQhOCq/+oub2oc5Ju/i/fd
iBWQL+N+gwxWUtVudDFMXheYG7iHjMXHbeEd2HyuOVSqY/9ytBRhSOE2UlbfErH0
Bvmgjj+Dg+e44nI4QnQxLhCFuVhtFS29fc9QYkaEuxleI0u5htoNHOvBmwDkhRmV
qJPJiyus/p5EVn5jzORxgG3Tf3xsiHAbI3TQzTRB4Cg/rxQ8mwHy2DxwJu8iFX77
hHWQpHNLh0gN/tUK7SWLnIPgYc98c2YMkv6Lmfj3OIEBj0IzmY3c1TqsyHXB54SS
+VXyeN0urYmxC3S8aTLglrtePr0faA1ytWh/qL/kU+yyEE+9I5cK8ablFk2yW1nZ
BOy+TEyDgdSkaBxTToa2N7ppQ92uuOxc68DP6+bP1QvkaD9iux1J3dgNivzBQ9tP
l+f3V8C6SLDkCAYQ+IVeqLpgfIRPi4IT568/BfZhQ9WFABwElXY9v4OM+BWfmk0J
4VLEO53rYLCF3j0bLoRZb1WH+x3jiwKnCe8bhIHAdzW84LAK8mwkYC0mw7NNM4Zt
wbA3XKPLicSK4vTk4e97n7GrYsREwxLau12wYWHRpPicLA78rD1ZXzPJgJAWDSX/
kbMBYrr/wFZQq8fNaN/zDgKQRyqTfKBSukO6yK53utb7dFbRQePhsMI9O7nIqv3c
Pe51nyLEFqfgj9Bmoy9NyinruhE1hSAEZ7FRWrki6YVH4eg93d08hAsLd8VaVtoP
32MUBRQO5RsseG6CyK9Pims7tMsOiQqNiVE31NrVDf44eveWoncK5GHXHqSlcS0Q
mZCo2WfUBDOWUYF4KRRLd5BQ1IevwK5ouVKDUi3Ek29d4heh6Gmls6VcMswwxOAi
0e8G5OSm4EE76uaBJmyBYupYB6PsJC4kFj7pbCweSRGKP9ESHjrRdei6SO8Wh3wg
1s/qgQczsbs270KXsS+8WcrSCDcTcmDTeEXT6oRXnaWtOoAT6Yc9on5009gU1rCT
hW6PdwaC5v0cCHR07C5M5QTOZxpAwqU6O+V01cjUlmkbYdHBG1epOOTEQhAr/ATe
ra/k0xUhqEoEqFVmEsZmIix7ZSl4z50jcLMCiDraqa74T5CpLX3HQB9HuNQcCmtf
WM/JPmJfgjQ6QfrhUSomfA48gqXRfhcTVM5E4CrEAEMVcRUFIhphBwr4ClJl347h
IpicwY8u+sFktrUfJfOazZwb0zHpO0UQ7nC/RHQGgQYr2c4TilnwZoDl4j12kATq
CwjCXVCDzf6reaFzKvNeozwEFkeTXrvdnu66UssoP18qokNEP5F2jJPU2MxzjAls
Se63knt3XLkumjFmF0YkrBCfqoBG7vGNkMK8KM+mPAGwOxZjHij0281k/uWcJc/x
3L9bYXyu/94AtL25UPxb/0VIGt9zZQO7G7hu32h2iqvemEFmwzRHkurqmeR6PgW/
5qWuk0WvebOo7R64HPlNiUi5L/Ik/CVz4Jje+NG3XtKHRW4jiFHS0GBwhE/lawWC
eKTAU6pxtBZ3Ws88w1GqSq8lKiP39QUpRuROWBmVrKF+mL/2eVKXmQ/0EJqwtFSf
dy0EZbp6RXk8+xW9bdtua2rgKZ4QzLfUz/tjfMNRbgZVFFvn3N/Yrz4UjcG+n2wA
Q5wzEfNrh6dM611tW+Ts7ioYsMP8RDoOX4ftBtpjJ6ecwSfTWCQkiacpgvojfB+N
/Pidx3U/Xt41IqG5a6k3QBFKTfCRc5SQLEZjl2UPo0XajyuuOEgnMBAV6Eqani2L
Xbr3PiW+4a3/VWUBc26jd3ZCaoSDhxhtUlZDLUlu0z+xHCszFiHpHO0BI2/bKiia
oNZlhYQjOO2QtKp9WbHfDWe/cIfzOrjU6Y4d/iNihVLldSqLRuoDknT3e+0vC9BV
B5s3DBJFm9rB3R6bsQdON1I/AgPmPnWNPf+cNV8yDOTNa9eJs+zc+xXZtgPoOXNm
Ud0d4MrUf5umxu8yUio90Sdva1R4jTqMP1iOh18k71ZJAg1JYDrptoxa9/y2DdnD
RxYuT6uoUAC01SYfBPjiwSgH1xtF3eP4IQBa5ZnWD7gK4enZwZXsowrQ+Vu0jcJ7
S945U89pKflXdfOi95DIvM2KRoljAJPN2ZEP1bjbfTRZA/wA4yxaeSijNA/U45FH
uOAHBM66U9oeLgX+MgcHlbDYVw9ig/rsvQeqfoLnQQOlqjQg5bHbqHlrUzAVE0FM
WcGnf/o/BpQGbcwqLOC1EPI3O6zTyJRFzrRw7g/rCx69aObNYhogSiOzYwd0MIqk
/fWD3N2uf7+UPE9PKede2GjnL6RlDvD4Jpxa9AziYb5gmfhyevrxFXXpjiKq8LIh
53AuVcnXV35DF1DwF1CsbvTpvZQNI9rJXRPiwfvQnKNj5UNUJXcHpqGA4ZqfLGPN
cpCCrYAhD47ZiEDSAeM7EuWVByXR88qLbeK49wCmPitFM/xxg34OhlnaLDO/hGa2
+Yuakonfcz8vn0kk5DMvuTbYuGgBWevPAkk1B0+oy9sYabAUUj+bdsnEoSclCtgJ
2Y3+8ziOIlDi5VR+gjnSTLwo52rvRDiovHfFBiWaWBrI63/WYpqdKs7Rmg3Fl6J9
J0k4tjw5TPAhVR87rvusTfwBjNPo4JmqKFgKUxYe1DFCpoALGZCaoS8hpTwBjrZ6
C1l7PAVsXN/XwBkV13FQl050XNuUk/yhAkpq3Pt3TadiubCoyLzX2jnojbDj3oUr
TX6ur0rU1CVyG2QZX+0/peXLcdLqmVrQb4ld/IlvCU1ZZwTcr8pxS7JKsaqQdT7y
reFP45kony/2sVSFHujA9tJIWvESJD6yWptdnGTuiaQZflyC444LxpPutULE8/nr
/byxnGToGV4ic5ftr/fMwvCEKHtNa6RA+1UmWESo4po7hba3zWETZees0YvV3KRC
lpjHor9X6XAxYpHgUweW1MUSJB8o+MSjPkfriR79JBYKMdwVDY9Fv07R9Er1fcuw
gp/G6JujqXw17UAHzh6CuCxQd2T6rDNmJe2QScvEMYoEhTpVyaExf85KuqrqgTU4
VGUxweD6fFM7IZclgOvno9pz35285U82JdNdlRCIfwH70AMBJKmkYsXb2hRtub7c
5/suDk6u8Khvaf3oEhKNURDgjIatYuP2/Ux9YzZfvTQQVccrCvTEqPnMjduQl+6o
kqM9LDI00dLm/vGJa4Ld2W/0AeQhNvFGxgcN0bCbp4t97UxIU9l3NIvnpFF2Zx+8
IMvQ1cytjxOqLD9KPGR1izXbd5MYn8JB3C2sjQreVQ7eVy36/NqQDEbcQegtuH6Y
t5HjwVcHUcSgKorGvZrAWRT4XXQtb79vLhxljry8758V7UwXAt/IF2IImQ9ZB8O9
ggJu/EJJIfqK8l7txXvocG0IZcn8E8mQu1GfkAn6IrB68euLYDIwUfa6xUeGbxZe
zqW0UeRyWx40sybd82vnZaS26MBG5X7pQ4400v7Nxhdp8KJ2wm4rX2BJsLzvIQeU
yM/rpGDzlzLGRmTLnV10HuCImVVJ6uvi10Jdx3O5lfxQZ+PT5GCEHL5WF30AXrnG
D16s36UdcJ+avF3XA/AmDW4aeHxu+JRSCvBDhQCiRQm1SFM8PfWOCFlXgPM9GA6P
RdiR5J6AiovalUagiKb0cvAqUSD0w1IYkmpd24XX1ax+iL9ACuvH9bhyJB3gvEyJ
gueYzT0VCz3ETZIFte7EV2oGTFiVrQ9mD4Jri1QShpo3kbhQgc4veIH40q9Unb4I
JALCqzhi0R3G9D7aLNaAN75c1E52Fw5Vv6yiNQ+VGg/IKZ50GP0jSlnw0IuZ4Qiw
`protect end_protected